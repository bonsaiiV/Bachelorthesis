library ieee;
use ieee.std_logic_1164.all;
entity fft_tb is
end fft_tb;
architecture test of fft_tb is
    component fft
    port (
       clk, fft_start: in std_logic;
       output_valid : out std_logic;
       inA, inB : in std_logic_vector(47 downto 0);
       outA, outB: out std_logic_vector(47 downto 0));
    end component;
signal inA, inB, outA, outB : std_logic_vector(47 downto 0) := (others =>'0');
    signal clk, fft_start : std_logic := '0';
    signal output_valid : std_logic;
begin
    fft_i: fft
    port map (
        clk => clk,
        fft_start => fft_start,
        inA => inA,
        inB => inB,
        output_valid => output_valid,
        outA => outA,
        outB => outB
    );
   process begin
        wait for 1 ns;
        clk <= '1';
        wait for 1 ns;
        clk <= '0';
        fft_start <= '1';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000100100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110001110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000100010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000111110101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101111110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000111110101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000100101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000100011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000101100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000110000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111110100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111110100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000101000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101111010000000000000";
inB<="000000000000000000000000000100000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000100110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000011111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111110010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111110100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100011010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000100000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111110100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000111110111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000111110111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100101110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111110011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000100011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100110010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111110111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101001000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111110111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000100001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000111110111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100111010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111110100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000100011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111101100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000011111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101000010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000011111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111110010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110000100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000100100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000011111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110000000000000000";
inB<="000000000000000000000000000100111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000100100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111110100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000111110101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111110001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000100001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110000000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111110000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111110101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111101110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111110111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000100110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100101000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000111101111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000100010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000101010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000100011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000011111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000100001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111110101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111110010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000100010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111110111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111110000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110000000000000000";
inB<="000000000000000000000000111110010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000111110100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000100111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000100001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111110010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010110000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000111110001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111100000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000100101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000100001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101001100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000100011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000011110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110001110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111101110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101011100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110000100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000100001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000011111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110000110000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000100010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000100101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111110000000000000";
inB<="000000000000000000000000000011111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111110101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100111100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111110110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111110110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111110110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111110101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110001100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000101000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000011110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101110010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000100011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000100101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000100110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111110100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100100000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000100010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101001110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111110010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111110010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111110111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000100000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000100010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000011111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100101100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100111000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000011110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000100010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000100010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000011110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011100000000000000";
inB<="000000000000000000000000000100011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111110100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101001010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000100111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111110100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000100100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100011110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000100101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111110101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101010000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111110100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001000000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000100001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000111110111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000101010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111110101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101101000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111110011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000100010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000100100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000100110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000011110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111110001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101111110000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000100001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000100010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000111110011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100011110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111110100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110001000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000100011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000111110101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000111110111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100111010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000100001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110001100000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110000000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000100000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111110011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000111110100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011010000000000000";
inB<="000000000000000000000000000100011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000111110111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000100010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000100000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000100001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000011110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000100100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000100001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000111110110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111110001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111101110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111110111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000100110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000100010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000011111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110000000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111110110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111110001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100101000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111110011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000011111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000101011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111110100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000100011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000011111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000100010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111100000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111110101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101000010000000000000";
inB<="000000000000000000000000111110001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101011010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111110001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100101100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100101010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101011110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100101100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000111110101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111110010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000011111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110000110000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111110111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000100101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000100110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111110011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010010000000000000";
inB<="000000000000000000000000111110010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000100001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111110111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101010100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111110101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111110100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011010000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111110100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111110100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000011111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000100000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000111110110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101000100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000100101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110001100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000100001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000100010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000111110001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000100110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111101011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111110101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010000000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111110100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000110010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000100011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111110111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000100100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111110101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111110010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000100001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100101110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101001010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111110111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000101011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000100001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101110010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000100011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100011010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111110010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000011111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000011111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010000000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100011010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000100010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100101010000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000100110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110001010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000011111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000111110011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111110100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111110111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000100010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111110101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000101000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101000100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101010000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101100100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000100110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111101111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111110000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000100011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111110100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101111110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000100111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000100011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110001110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110001000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000100000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111101000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000100000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111110000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101101000000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000111110100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111110100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111110000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100111000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000111110111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101010010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000101000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100011010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000111110101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000100101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111110101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101110110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100011010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000111110000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101010000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000100001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111101111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000100110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100011010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000100000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000111110100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110000010000000000000";
inB<="000000000000000000000000000101101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000100000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101111000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111100110110000000000000";
inB<="000000000000000000000000000100001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101101010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111110111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111110111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000111101111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000011110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111110000000000000";
inB<="000000000000000000000000111101111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100110010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100110000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011100000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000100001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111110111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000100010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000111110101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000100110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000100101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111110100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111100000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000100001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000100000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111110111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100011110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000100011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100011110000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100111000000000000000";
inB<="000000000000000000000000111110111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111110111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000111110100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100000000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111101110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111110111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000100010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101001000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110001000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101011000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111110110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111101000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111010000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110000010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000100100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000101000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000100010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000011111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000111110010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000100001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100110010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100011000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111110011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000111110101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000100101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000011111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111110111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100101000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000100011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000100000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110010000000000000";
inB<="000000000000000000000000000100100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101001000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000100110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000011110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101100100000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000100101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000111110110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111110100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000101011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100110010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111110011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000100010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111110100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101110010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000111110100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000100111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000100000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000111110100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110001110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000111110111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000111110010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111110011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000111110111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111110101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100101100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000100101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000100100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011110000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111110000000000000";
inB<="000000000000000000000000111110100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111110001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111110011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100111100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000100001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110001100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101111000000000000000";
inB<="000000000000000000000000111110101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111110011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000100000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000100010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000100000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100011110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000111110111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000100000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000100000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000100010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100110000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111110011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111110110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111110111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000101001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010110000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111110010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000100111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000100101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000111110110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000100101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000100001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111110011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111110000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110001110000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110000000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100010000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000100001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000100000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000111110100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111110001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000100010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000110000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000011111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000100011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111110011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111101111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111000000000000000";
inB<="000000000000000000000000000100101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001010000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000111110110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000111101111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100000000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101100010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111110011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000100000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000100000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110010000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111110111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111110110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101010010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000111101110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000011111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111100110000000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000100110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101101010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110100110000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000100011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000100000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111101101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000100010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100101110000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000011101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111110010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101000000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000111110111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000100001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101011010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000011100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000100101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100110110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000101000000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111100000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100010000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111000110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000011100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000100100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000100010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111110110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000100011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000110000000000000";
inB<="000000000000000000000000111111001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101110100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111010000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000011111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000011010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000111111000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111110011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100010000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000011011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000100011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000100001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000011110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000100000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000100000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101010000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000111110111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100001100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000100101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000011000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011111000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000111110101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110010000000000000";
inB<="000000000000000000000000000011110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111110110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000011100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000011000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010000000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110110000000000000";
inB<="000000000000000000000000111111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000111111001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000100000000000000";
inB<="000000000000000000000000000011001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000111111001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001010000000000000";
inB<="000000000000000000000000000101000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110111010000000000000";
inB<="000000000000000000000000111111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000011000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011000000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010000000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000011100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000010000000000000";
inB<="000000000000000000000000000010101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010100000000000000";
inB<="000000000000000000000000000010100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000100110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000001010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000011101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111100000000000000";
inB<="000000000000000000000000000011111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000111110111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001100000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000111111000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000111110010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000100000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111101101000000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011010000000000000";
inB<="000000000000000000000000111111000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000011010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000011010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000011110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110100000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000011011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101010000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011010000000000000";
inB<="000000000000000000000000111110100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001110000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000111110110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100000000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000111111010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000010111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111110000000000000";
inB<="000000000000000000000000000011010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111110111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010110000000000000";
inB<="000000000000000000000000000010111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110110110000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010010000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110110000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001010000000000000";
inB<="000000000000000000000000000000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110110000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000100000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000111110111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000100001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110000000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000111111010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000000011001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000000000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000111111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011001000000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000011101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000001101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110010110000000000000";
inB<="000000000000000000000000000001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111100000000000000";
inB<="000000000000000000000000000011001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110101100000000000000";
inB<="000000000000000000000000000001111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111000000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100010000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000110000000000000";
inB<="000000000000000000000000000010100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000001110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100000000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111111010000000000000";
inB<="000000000000000000000000000011000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000111111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000110000000000000";
inB<="000000000000000000000000000001101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011110000000000000";
inB<="000000000000000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001010000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100110000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000010010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100100100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011110010000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110010000000000000";
inB<="000000000000000000000000000001101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000100000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000111111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000010101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010100000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000000000000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011000000000000000";
inB<="000000000000000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000010000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101000000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110100000000000000";
inB<="000000000000000000000000000010110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101100000000000000";
inB<="000000000000000000000000000010101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000111111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010000000000000000";
inB<="000000000000000000000000000010110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111110011100000000000000";
inB<="000000000000000000000000000011111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011100000000000000";
inB<="000000000000000000000000000000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011100110000000000000";
inB<="000000000000000000000000000000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000010000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111100100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101110000000000000";
inB<="000000000000000000000000000010011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111010000000000000";
inB<="000000000000000000000000000011011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000000001100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011010110000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001000000000000000";
inB<="000000000000000000000000000010011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111110000000000000000";
inB<="000000000000000000000000000000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101000000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111110000000000000";
inB<="000000000000000000000000000001100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110100000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111011110000000000000";
inB<="000000000000000000000000111111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111010110000000000000";
inB<="000000000000000000000000000100111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011110000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000111111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100010000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011000000000000000";
inB<="000000000000000000000000000010011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000000000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000000000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010110000000000000";
inB<="000000000000000000000000000010100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000010110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000110100000000000000";
inB<="000000000000000000000000000001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000100110000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000001111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001000000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010010000000000000";
inB<="000000000000000000000000000001101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110110000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111110000000000000";
inB<="000000000000000000000000000001001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011011100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000000000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001100000000000000";
inB<="000000000000000000000000000001100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111010000000000000";
inB<="000000000000000000000000000000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000111111001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101000000000000000";
inB<="000000000000000000000000000010010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000111111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000100000000000000000000";
inB<="000000000000000000000000111111011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010110000000000000";
inB<="000000000000000000000000000010001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001010000000000000";
inB<="000000000000000000000000000001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000011100000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000010011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000011101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111100000000000000";
inB<="000000000000000000000000000001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111101110000000000000";
inB<="000000000000000000000000111110111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010100110000000000000";
inB<="000000000000000000000000000010001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000001110000000000000";
inB<="000000000000000000000000111110010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101010000000000000";
inB<="000000000000000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101100000000000000";
inB<="000000000000000000000000000001110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011100000000000000";
inB<="000000000000000000000000000010001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101000000000000000";
inB<="000000000000000000000000111111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001110010000000000000";
inB<="000000000000000000000000000000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001100110000000000000";
inB<="000000000000000000000000000000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010000000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000100000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010010100000000000000";
inB<="000000000000000000000000000001100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010100000000000000";
inB<="000000000000000000000000111111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010110000000000000000";
inB<="000000000000000000000000000000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001100000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000111000000000000000";
inB<="000000000000000000000000000001011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000111111001000000000000000";
inB<="000000000000000000000000000010010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000010010000000000000";
inB<="000000000000000000000000000001110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001000000000000000";
inB<="000000000000000000000000000000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001101110000000000000";
inB<="000000000000000000000000000010100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001100000000000000";
inB<="000000000000000000000000111111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111110000000000000";
inB<="000000000000000000000000000000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101010000000000000";
inB<="000000000000000000000000000001011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111110111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011101110000000000000";
inB<="000000000000000000000000000010000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001011000000000000000";
inB<="000000000000000000000000111111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010000000000000000000";
inB<="000000000000000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001000000000000000000";
inB<="000000000000000000000000111111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010111010000000000000";
inB<="000000000000000000000000111111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010011110000000000000";
inB<="000000000000000000000000111111010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001010010000000000000";
inB<="000000000000000000000000000000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000011000110000000000000";
inB<="000000000000000000000000000000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010101100000000000000";
inB<="000000000000000000000000000000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001111000000000000000";
inB<="000000000000000000000000000000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000010001010000000000000";
inB<="000000000000000000000000000001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000000101110000000000000";
inB<="000000000000000000000000000011001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000000001001110000000000000";
inB<="000000000000000000000000000001101010000000000000";
while output_valid = '0' loop
            wait for 1 ns;
            clk <= '1';
            wait for 1 ns;
            clk <= '0';
        end loop;
        for i in 0 to 16384 loop
        wait for 1 ns;
            clk <= '1';
            wait for 1 ns;
            clk <= '0';
        end loop;
        wait;
    end process;
end test;
