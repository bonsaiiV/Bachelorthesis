library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity rom is
    generic(
        width :integer:=12;
        length :integer
    ) ;
    port (
       clk: std_logic;
       addr: in std_logic_vector(length-1 downto 0);
       value: out std_logic_vector(width-1 downto 0)
    );
end rom;
architecture rom_b of rom is
    type MEMORY is array(0 to 2**length-1) of std_logic_vector(width-1 downto 0);
    signal rom_mem :MEMORY :=(
"00000000000100000000","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","00000000000011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111110011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111100011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111010011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111111000011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110110011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110100011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110010011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111110000011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101110011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101100011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101010011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111101000011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100110011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100100011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100010011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111100000011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011110011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011100011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011010011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111011000011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010110011111111","11111010100011111111","11111010100011111111","11111010100011111111","11111010100011111111","11111010100011111111","11111010100011111111","11111010100011111111","11111010100011111111","11111010100011111111","11111010100011111111","11111010100011111111","11111010100011111111","11111010100011111111","11111010100011111110","11111010100011111110","11111010100011111110","11111010100011111110","11111010100011111110","11111010100011111110","11111010100011111110","11111010100011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010010011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111010000011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001110011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001100011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001010011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111001000011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000110011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000100011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111110","11111000010011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11111000000011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111110011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111100011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111010011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110111000011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110110011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110100011111101","11110110010011111101","11110110010011111101","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110010011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110110000011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101110011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101100011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101010011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110101000011111100","11110100110011111100","11110100110011111100","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100110011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100100011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100010011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110100000011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011110011111011","11110011100011111011","11110011100011111011","11110011100011111011","11110011100011111011","11110011100011111011","11110011100011111011","11110011100011111011","11110011100011111010","11110011100011111010","11110011100011111010","11110011100011111010","11110011100011111010","11110011100011111010","11110011100011111010","11110011100011111010","11110011100011111010","11110011100011111010","11110011100011111010","11110011100011111010","11110011100011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011010011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110011000011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010110011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010100011111010","11110010010011111010","11110010010011111010","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010010011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110010000011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001110011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001100011111001","11110001010011111001","11110001010011111001","11110001010011111001","11110001010011111001","11110001010011111001","11110001010011111001","11110001010011111001","11110001010011111001","11110001010011111001","11110001010011111001","11110001010011111000","11110001010011111000","11110001010011111000","11110001010011111000","11110001010011111000","11110001010011111000","11110001010011111000","11110001010011111000","11110001010011111000","11110001010011111000","11110001010011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110001000011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000110011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000100011111000","11110000010011111000","11110000010011111000","11110000010011111000","11110000010011111000","11110000010011111000","11110000010011111000","11110000010011111000","11110000010011111000","11110000010011111000","11110000010011111000","11110000010011111000","11110000010011110111","11110000010011110111","11110000010011110111","11110000010011110111","11110000010011110111","11110000010011110111","11110000010011110111","11110000010011110111","11110000010011110111","11110000010011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11110000000011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111110011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111100011110111","11101111010011110111","11101111010011110111","11101111010011110111","11101111010011110111","11101111010011110111","11101111010011110111","11101111010011110110","11101111010011110110","11101111010011110110","11101111010011110110","11101111010011110110","11101111010011110110","11101111010011110110","11101111010011110110","11101111010011110110","11101111010011110110","11101111010011110110","11101111010011110110","11101111010011110110","11101111010011110110","11101111010011110110","11101111010011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101111000011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110110011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110110","11101110100011110101","11101110100011110101","11101110100011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110010011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101110000011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101110011110101","11101101100011110101","11101101100011110101","11101101100011110101","11101101100011110101","11101101100011110101","11101101100011110100","11101101100011110100","11101101100011110100","11101101100011110100","11101101100011110100","11101101100011110100","11101101100011110100","11101101100011110100","11101101100011110100","11101101100011110100","11101101100011110100","11101101100011110100","11101101100011110100","11101101100011110100","11101101100011110100","11101101100011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101010011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101101000011110100","11101100110011110100","11101100110011110100","11101100110011110100","11101100110011110100","11101100110011110100","11101100110011110100","11101100110011110100","11101100110011110100","11101100110011110100","11101100110011110100","11101100110011110011","11101100110011110011","11101100110011110011","11101100110011110011","11101100110011110011","11101100110011110011","11101100110011110011","11101100110011110011","11101100110011110011","11101100110011110011","11101100110011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100100011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100010011110011","11101100000011110011","11101100000011110011","11101100000011110011","11101100000011110011","11101100000011110011","11101100000011110011","11101100000011110011","11101100000011110011","11101100000011110011","11101100000011110011","11101100000011110011","11101100000011110011","11101100000011110010","11101100000011110010","11101100000011110010","11101100000011110010","11101100000011110010","11101100000011110010","11101100000011110010","11101100000011110010","11101100000011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011110011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011100011110010","11101011010011110010","11101011010011110010","11101011010011110010","11101011010011110010","11101011010011110010","11101011010011110010","11101011010011110010","11101011010011110010","11101011010011110010","11101011010011110010","11101011010011110010","11101011010011110001","11101011010011110001","11101011010011110001","11101011010011110001","11101011010011110001","11101011010011110001","11101011010011110001","11101011010011110001","11101011010011110001","11101011010011110001","11101011010011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101011000011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010110011110001","11101010100011110001","11101010100011110001","11101010100011110001","11101010100011110001","11101010100011110001","11101010100011110001","11101010100011110001","11101010100011110001","11101010100011110000","11101010100011110000","11101010100011110000","11101010100011110000","11101010100011110000","11101010100011110000","11101010100011110000","11101010100011110000","11101010100011110000","11101010100011110000","11101010100011110000","11101010100011110000","11101010100011110000","11101010100011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010010011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101010000011110000","11101001110011110000","11101001110011110000","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001110011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001100011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101111","11101001010011101110","11101001010011101110","11101001010011101110","11101001010011101110","11101001010011101110","11101001010011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101001000011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000110011101110","11101000100011101110","11101000100011101110","11101000100011101110","11101000100011101110","11101000100011101110","11101000100011101110","11101000100011101110","11101000100011101101","11101000100011101101","11101000100011101101","11101000100011101101","11101000100011101101","11101000100011101101","11101000100011101101","11101000100011101101","11101000100011101101","11101000100011101101","11101000100011101101","11101000100011101101","11101000100011101101","11101000100011101101","11101000100011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000010011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101101","11101000000011101100","11101000000011101100","11101000000011101100","11101000000011101100","11101000000011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111110011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111100011101100","11100111010011101100","11100111010011101100","11100111010011101100","11100111010011101100","11100111010011101100","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111010011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100111000011101011","11100110110011101011","11100110110011101011","11100110110011101011","11100110110011101011","11100110110011101011","11100110110011101011","11100110110011101011","11100110110011101011","11100110110011101011","11100110110011101011","11100110110011101011","11100110110011101011","11100110110011101010","11100110110011101010","11100110110011101010","11100110110011101010","11100110110011101010","11100110110011101010","11100110110011101010","11100110110011101010","11100110110011101010","11100110110011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110100011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101010","11100110010011101001","11100110010011101001","11100110010011101001","11100110010011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100110000011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101110011101001","11100101100011101001","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101100011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101010011101000","11100101000011101000","11100101000011101000","11100101000011101000","11100101000011101000","11100101000011101000","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100101000011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100110011100111","11100100100011100111","11100100100011100111","11100100100011100111","11100100100011100111","11100100100011100111","11100100100011100111","11100100100011100111","11100100100011100110","11100100100011100110","11100100100011100110","11100100100011100110","11100100100011100110","11100100100011100110","11100100100011100110","11100100100011100110","11100100100011100110","11100100100011100110","11100100100011100110","11100100100011100110","11100100100011100110","11100100100011100110","11100100100011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100010011100110","11100100000011100110","11100100000011100110","11100100000011100110","11100100000011100110","11100100000011100110","11100100000011100110","11100100000011100110","11100100000011100110","11100100000011100110","11100100000011100101","11100100000011100101","11100100000011100101","11100100000011100101","11100100000011100101","11100100000011100101","11100100000011100101","11100100000011100101","11100100000011100101","11100100000011100101","11100100000011100101","11100100000011100101","11100100000011100101","11100100000011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011110011100101","11100011100011100101","11100011100011100101","11100011100011100101","11100011100011100101","11100011100011100101","11100011100011100101","11100011100011100101","11100011100011100101","11100011100011100101","11100011100011100101","11100011100011100100","11100011100011100100","11100011100011100100","11100011100011100100","11100011100011100100","11100011100011100100","11100011100011100100","11100011100011100100","11100011100011100100","11100011100011100100","11100011100011100100","11100011100011100100","11100011100011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011010011100100","11100011000011100100","11100011000011100100","11100011000011100100","11100011000011100100","11100011000011100100","11100011000011100100","11100011000011100100","11100011000011100100","11100011000011100100","11100011000011100011","11100011000011100011","11100011000011100011","11100011000011100011","11100011000011100011","11100011000011100011","11100011000011100011","11100011000011100011","11100011000011100011","11100011000011100011","11100011000011100011","11100011000011100011","11100011000011100011","11100011000011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010110011100011","11100010100011100011","11100010100011100011","11100010100011100011","11100010100011100011","11100010100011100011","11100010100011100011","11100010100011100011","11100010100011100011","11100010100011100010","11100010100011100010","11100010100011100010","11100010100011100010","11100010100011100010","11100010100011100010","11100010100011100010","11100010100011100010","11100010100011100010","11100010100011100010","11100010100011100010","11100010100011100010","11100010100011100010","11100010100011100010","11100010100011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010010011100010","11100010000011100010","11100010000011100010","11100010000011100010","11100010000011100010","11100010000011100010","11100010000011100010","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100010000011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001110011100001","11100001100011100001","11100001100011100001","11100001100011100001","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001100011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011100000","11100001010011011111","11100001010011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100001000011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011111","11100000110011011110","11100000110011011110","11100000110011011110","11100000110011011110","11100000110011011110","11100000110011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000100011011110","11100000010011011110","11100000010011011110","11100000010011011110","11100000010011011110","11100000010011011110","11100000010011011110","11100000010011011110","11100000010011011110","11100000010011011110","11100000010011011110","11100000010011011110","11100000010011011101","11100000010011011101","11100000010011011101","11100000010011011101","11100000010011011101","11100000010011011101","11100000010011011101","11100000010011011101","11100000010011011101","11100000010011011101","11100000010011011101","11100000010011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11100000000011011101","11011111110011011101","11011111110011011101","11011111110011011101","11011111110011011101","11011111110011011101","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111110011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011100","11011111100011011011","11011111100011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111010011011011","11011111000011011011","11011111000011011011","11011111000011011011","11011111000011011011","11011111000011011011","11011111000011011011","11011111000011011011","11011111000011011011","11011111000011011011","11011111000011011011","11011111000011011011","11011111000011011011","11011111000011011011","11011111000011011010","11011111000011011010","11011111000011011010","11011111000011011010","11011111000011011010","11011111000011011010","11011111000011011010","11011111000011011010","11011111000011011010","11011111000011011010","11011111000011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110110011011010","11011110100011011010","11011110100011011010","11011110100011011010","11011110100011011010","11011110100011011010","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110100011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011001","11011110010011011000","11011110010011011000","11011110010011011000","11011110010011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011110000011011000","11011101110011011000","11011101110011011000","11011101110011011000","11011101110011011000","11011101110011011000","11011101110011011000","11011101110011011000","11011101110011011000","11011101110011011000","11011101110011011000","11011101110011010111","11011101110011010111","11011101110011010111","11011101110011010111","11011101110011010111","11011101110011010111","11011101110011010111","11011101110011010111","11011101110011010111","11011101110011010111","11011101110011010111","11011101110011010111","11011101110011010111","11011101110011010111","11011101110011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010111","11011101100011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101010011010110","11011101000011010110","11011101000011010110","11011101000011010110","11011101000011010110","11011101000011010110","11011101000011010110","11011101000011010110","11011101000011010110","11011101000011010110","11011101000011010110","11011101000011010110","11011101000011010110","11011101000011010101","11011101000011010101","11011101000011010101","11011101000011010101","11011101000011010101","11011101000011010101","11011101000011010101","11011101000011010101","11011101000011010101","11011101000011010101","11011101000011010101","11011101000011010101","11011101000011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100110011010101","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100100011010100","11011100010011010100","11011100010011010100","11011100010011010100","11011100010011010100","11011100010011010100","11011100010011010100","11011100010011010100","11011100010011010100","11011100010011010100","11011100010011010100","11011100010011010100","11011100010011010100","11011100010011010100","11011100010011010011","11011100010011010011","11011100010011010011","11011100010011010011","11011100010011010011","11011100010011010011","11011100010011010011","11011100010011010011","11011100010011010011","11011100010011010011","11011100010011010011","11011100010011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010011","11011100000011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011110011010010","11011011100011010010","11011011100011010010","11011011100011010010","11011011100011010010","11011011100011010010","11011011100011010010","11011011100011010010","11011011100011010010","11011011100011010010","11011011100011010010","11011011100011010001","11011011100011010001","11011011100011010001","11011011100011010001","11011011100011010001","11011011100011010001","11011011100011010001","11011011100011010001","11011011100011010001","11011011100011010001","11011011100011010001","11011011100011010001","11011011100011010001","11011011100011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010001","11011011010011010000","11011011010011010000","11011011010011010000","11011011010011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011011000011010000","11011010110011010000","11011010110011010000","11011010110011010000","11011010110011010000","11011010110011010000","11011010110011010000","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010110011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001111","11011010100011001110","11011010100011001110","11011010100011001110","11011010100011001110","11011010100011001110","11011010100011001110","11011010100011001110","11011010100011001110","11011010100011001110","11011010100011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010010011001110","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011010000011001101","11011001110011001101","11011001110011001101","11011001110011001101","11011001110011001101","11011001110011001101","11011001110011001101","11011001110011001101","11011001110011001101","11011001110011001101","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001110011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001100","11011001100011001011","11011001100011001011","11011001100011001011","11011001100011001011","11011001100011001011","11011001100011001011","11011001100011001011","11011001100011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001011","11011001010011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011001000011001010","11011000110011001010","11011000110011001010","11011000110011001010","11011000110011001010","11011000110011001010","11011000110011001010","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000110011001001","11011000100011001001","11011000100011001001","11011000100011001001","11011000100011001001","11011000100011001001","11011000100011001001","11011000100011001001","11011000100011001001","11011000100011001001","11011000100011001001","11011000100011001001","11011000100011001001","11011000100011001001","11011000100011001001","11011000100011001000","11011000100011001000","11011000100011001000","11011000100011001000","11011000100011001000","11011000100011001000","11011000100011001000","11011000100011001000","11011000100011001000","11011000100011001000","11011000100011001000","11011000100011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011001000","11011000010011000111","11011000010011000111","11011000010011000111","11011000010011000111","11011000010011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11011000000011000111","11010111110011000111","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111110011000110","11010111100011000110","11010111100011000110","11010111100011000110","11010111100011000110","11010111100011000110","11010111100011000110","11010111100011000110","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111100011000101","11010111010011000101","11010111010011000101","11010111010011000101","11010111010011000101","11010111010011000101","11010111010011000101","11010111010011000101","11010111010011000101","11010111010011000101","11010111010011000101","11010111010011000101","11010111010011000101","11010111010011000101","11010111010011000100","11010111010011000100","11010111010011000100","11010111010011000100","11010111010011000100","11010111010011000100","11010111010011000100","11010111010011000100","11010111010011000100","11010111010011000100","11010111010011000100","11010111010011000100","11010111010011000100","11010111010011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000100","11010111000011000011","11010111000011000011","11010111000011000011","11010111000011000011","11010111000011000011","11010111000011000011","11010111000011000011","11010111000011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000011","11010110110011000010","11010110110011000010","11010110110011000010","11010110110011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110100011000010","11010110010011000010","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110010011000001","11010110000011000001","11010110000011000001","11010110000011000001","11010110000011000001","11010110000011000001","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010110000011000000","11010101110011000000","11010101110011000000","11010101110011000000","11010101110011000000","11010101110011000000","11010101110011000000","11010101110011000000","11010101110011000000","11010101110011000000","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101110010111111","11010101100010111111","11010101100010111111","11010101100010111111","11010101100010111111","11010101100010111111","11010101100010111111","11010101100010111111","11010101100010111111","11010101100010111111","11010101100010111111","11010101100010111111","11010101100010111111","11010101100010111110","11010101100010111110","11010101100010111110","11010101100010111110","11010101100010111110","11010101100010111110","11010101100010111110","11010101100010111110","11010101100010111110","11010101100010111110","11010101100010111110","11010101100010111110","11010101100010111110","11010101100010111110","11010101100010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111110","11010101010010111101","11010101010010111101","11010101010010111101","11010101010010111101","11010101010010111101","11010101010010111101","11010101010010111101","11010101010010111101","11010101010010111101","11010101010010111101","11010101010010111101","11010101010010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111101","11010101000010111100","11010101000010111100","11010101000010111100","11010101000010111100","11010101000010111100","11010101000010111100","11010101000010111100","11010101000010111100","11010101000010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111100","11010100110010111011","11010100110010111011","11010100110010111011","11010100110010111011","11010100110010111011","11010100110010111011","11010100110010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111011","11010100100010111010","11010100100010111010","11010100100010111010","11010100100010111010","11010100100010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111010","11010100010010111001","11010100010010111001","11010100010010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111001","11010100000010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011110010111000","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011100010110111","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011010010110110","11010011000010110110","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010011000010110101","11010010110010110101","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010110010110100","11010010100010110100","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010100010110011","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010010010110010","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110001","11010010000010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010110000","11010001110010101111","11010001110010101111","11010001110010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101111","11010001100010101110","11010001100010101110","11010001100010101110","11010001100010101110","11010001100010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101110","11010001010010101101","11010001010010101101","11010001010010101101","11010001010010101101","11010001010010101101","11010001010010101101","11010001010010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101101","11010001000010101100","11010001000010101100","11010001000010101100","11010001000010101100","11010001000010101100","11010001000010101100","11010001000010101100","11010001000010101100","11010001000010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101100","11010000110010101011","11010000110010101011","11010000110010101011","11010000110010101011","11010000110010101011","11010000110010101011","11010000110010101011","11010000110010101011","11010000110010101011","11010000110010101011","11010000110010101011","11010000110010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101011","11010000100010101010","11010000100010101010","11010000100010101010","11010000100010101010","11010000100010101010","11010000100010101010","11010000100010101010","11010000100010101010","11010000100010101010","11010000100010101010","11010000100010101010","11010000100010101010","11010000100010101010","11010000100010101010","11010000100010101010","11010000010010101010","11010000010010101010","11010000010010101010","11010000010010101010","11010000010010101010","11010000010010101010","11010000010010101010","11010000010010101010","11010000010010101010","11010000010010101010","11010000010010101010","11010000010010101010","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000010010101001","11010000000010101001","11010000000010101001","11010000000010101001","11010000000010101001","11010000000010101001","11010000000010101001","11010000000010101001","11010000000010101001","11010000000010101001","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11010000000010101000","11001111110010101000","11001111110010101000","11001111110010101000","11001111110010101000","11001111110010101000","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111110010100111","11001111100010100111","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100110","11001111100010100101","11001111100010100101","11001111100010100101","11001111100010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100101","11001111010010100100","11001111010010100100","11001111010010100100","11001111010010100100","11001111010010100100","11001111010010100100","11001111010010100100","11001111010010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100100","11001111000010100011","11001111000010100011","11001111000010100011","11001111000010100011","11001111000010100011","11001111000010100011","11001111000010100011","11001111000010100011","11001111000010100011","11001111000010100011","11001111000010100011","11001111000010100011","11001111000010100011","11001111000010100011","11001110110010100011","11001110110010100011","11001110110010100011","11001110110010100011","11001110110010100011","11001110110010100011","11001110110010100011","11001110110010100011","11001110110010100011","11001110110010100011","11001110110010100011","11001110110010100011","11001110110010100011","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110110010100010","11001110100010100010","11001110100010100010","11001110100010100010","11001110100010100010","11001110100010100010","11001110100010100010","11001110100010100010","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110100010100001","11001110010010100001","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010100000","11001110010010011111","11001110010010011111","11001110010010011111","11001110010010011111","11001110010010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011111","11001110000010011110","11001110000010011110","11001110000010011110","11001110000010011110","11001110000010011110","11001110000010011110","11001110000010011110","11001110000010011110","11001110000010011110","11001110000010011110","11001110000010011110","11001110000010011110","11001101110010011110","11001101110010011110","11001101110010011110","11001101110010011110","11001101110010011110","11001101110010011110","11001101110010011110","11001101110010011110","11001101110010011110","11001101110010011110","11001101110010011110","11001101110010011110","11001101110010011110","11001101110010011110","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101110010011101","11001101100010011101","11001101100010011101","11001101100010011101","11001101100010011101","11001101100010011101","11001101100010011101","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011100","11001101100010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011011","11001101010010011010","11001101010010011010","11001101010010011010","11001101010010011010","11001101010010011010","11001101010010011010","11001101010010011010","11001101010010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011010","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001101000010011001","11001100110010011001","11001100110010011001","11001100110010011001","11001100110010011001","11001100110010011001","11001100110010011001","11001100110010011001","11001100110010011001","11001100110010011001","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100110010011000","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010111","11001100100010010110","11001100100010010110","11001100100010010110","11001100100010010110","11001100100010010110","11001100100010010110","11001100100010010110","11001100100010010110","11001100100010010110","11001100100010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010110","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100010010010101","11001100000010010101","11001100000010010101","11001100000010010101","11001100000010010101","11001100000010010101","11001100000010010101","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010100","11001100000010010011","11001100000010010011","11001100000010010011","11001100000010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010011","11001011110010010010","11001011110010010010","11001011110010010010","11001011110010010010","11001011110010010010","11001011110010010010","11001011110010010010","11001011110010010010","11001011110010010010","11001011110010010010","11001011110010010010","11001011110010010010","11001011110010010010","11001011110010010010","11001011100010010010","11001011100010010010","11001011100010010010","11001011100010010010","11001011100010010010","11001011100010010010","11001011100010010010","11001011100010010010","11001011100010010010","11001011100010010010","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010001","11001011100010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010010000","11001011010010001111","11001011010010001111","11001011010010001111","11001011010010001111","11001011010010001111","11001011010010001111","11001011010010001111","11001011010010001111","11001011010010001111","11001011010010001111","11001011010010001111","11001011010010001111","11001011000010001111","11001011000010001111","11001011000010001111","11001011000010001111","11001011000010001111","11001011000010001111","11001011000010001111","11001011000010001111","11001011000010001111","11001011000010001111","11001011000010001111","11001011000010001111","11001011000010001111","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001011000010001110","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001101","11001010110010001100","11001010110010001100","11001010110010001100","11001010110010001100","11001010110010001100","11001010110010001100","11001010110010001100","11001010110010001100","11001010110010001100","11001010110010001100","11001010110010001100","11001010110010001100","11001010110010001100","11001010100010001100","11001010100010001100","11001010100010001100","11001010100010001100","11001010100010001100","11001010100010001100","11001010100010001100","11001010100010001100","11001010100010001100","11001010100010001100","11001010100010001100","11001010100010001100","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001011","11001010100010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001010","11001010010010001001","11001010010010001001","11001010010010001001","11001010010010001001","11001010010010001001","11001010010010001001","11001010010010001001","11001010010010001001","11001010010010001001","11001010010010001001","11001010010010001001","11001010010010001001","11001010010010001001","11001010010010001001","11001010010010001001","11001010000010001001","11001010000010001001","11001010000010001001","11001010000010001001","11001010000010001001","11001010000010001001","11001010000010001001","11001010000010001001","11001010000010001001","11001010000010001001","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010001000","11001010000010000111","11001010000010000111","11001010000010000111","11001010000010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000111","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001110010000110","11001001100010000110","11001001100010000110","11001001100010000110","11001001100010000110","11001001100010000110","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000101","11001001100010000100","11001001100010000100","11001001100010000100","11001001100010000100","11001001100010000100","11001001100010000100","11001001100010000100","11001001100010000100","11001001100010000100","11001001100010000100","11001001100010000100","11001001010010000100","11001001010010000100","11001001010010000100","11001001010010000100","11001001010010000100","11001001010010000100","11001001010010000100","11001001010010000100","11001001010010000100","11001001010010000100","11001001010010000100","11001001010010000100","11001001010010000100","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000011","11001001010010000010","11001001010010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000010","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001001000010000001","11001000110010000001","11001000110010000001","11001000110010000001","11001000110010000001","11001000110010000001","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110010000000","11001000110001111111","11001000110001111111","11001000110001111111","11001000110001111111","11001000110001111111","11001000110001111111","11001000110001111111","11001000110001111111","11001000110001111111","11001000110001111111","11001000110001111111","11001000110001111111","11001000100001111111","11001000100001111111","11001000100001111111","11001000100001111111","11001000100001111111","11001000100001111111","11001000100001111111","11001000100001111111","11001000100001111111","11001000100001111111","11001000100001111111","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111110","11001000100001111101","11001000100001111101","11001000100001111101","11001000100001111101","11001000100001111101","11001000100001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111101","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111100","11001000010001111011","11001000010001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111011","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11001000000001111010","11000111110001111010","11000111110001111010","11000111110001111010","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111001","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111110001111000","11000111100001111000","11000111100001111000","11000111100001111000","11000111100001111000","11000111100001111000","11000111100001111000","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110111","11000111100001110110","11000111100001110110","11000111100001110110","11000111100001110110","11000111100001110110","11000111100001110110","11000111100001110110","11000111100001110110","11000111100001110110","11000111100001110110","11000111100001110110","11000111100001110110","11000111100001110110","11000111100001110110","11000111100001110110","11000111010001110110","11000111010001110110","11000111010001110110","11000111010001110110","11000111010001110110","11000111010001110110","11000111010001110110","11000111010001110110","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110101","11000111010001110100","11000111010001110100","11000111010001110100","11000111010001110100","11000111010001110100","11000111010001110100","11000111010001110100","11000111010001110100","11000111010001110100","11000111010001110100","11000111010001110100","11000111010001110100","11000111010001110100","11000111010001110100","11000111000001110100","11000111000001110100","11000111000001110100","11000111000001110100","11000111000001110100","11000111000001110100","11000111000001110100","11000111000001110100","11000111000001110100","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110011","11000111000001110010","11000111000001110010","11000111000001110010","11000111000001110010","11000111000001110010","11000111000001110010","11000111000001110010","11000111000001110010","11000111000001110010","11000111000001110010","11000111000001110010","11000111000001110010","11000111000001110010","11000110110001110010","11000110110001110010","11000110110001110010","11000110110001110010","11000110110001110010","11000110110001110010","11000110110001110010","11000110110001110010","11000110110001110010","11000110110001110010","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110001","11000110110001110000","11000110110001110000","11000110110001110000","11000110110001110000","11000110110001110000","11000110110001110000","11000110110001110000","11000110110001110000","11000110110001110000","11000110110001110000","11000110110001110000","11000110110001110000","11000110110001110000","11000110110001110000","11000110100001110000","11000110100001110000","11000110100001110000","11000110100001110000","11000110100001110000","11000110100001110000","11000110100001110000","11000110100001110000","11000110100001110000","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101111","11000110100001101110","11000110100001101110","11000110100001101110","11000110100001101110","11000110100001101110","11000110100001101110","11000110100001101110","11000110100001101110","11000110100001101110","11000110100001101110","11000110100001101110","11000110100001101110","11000110100001101110","11000110100001101110","11000110100001101110","11000110010001101110","11000110010001101110","11000110010001101110","11000110010001101110","11000110010001101110","11000110010001101110","11000110010001101110","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101101","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110010001101100","11000110000001101100","11000110000001101100","11000110000001101100","11000110000001101100","11000110000001101100","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101011","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000110000001101010","11000101110001101010","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101001","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001101000","11000101110001100111","11000101110001100111","11000101110001100111","11000101110001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100111","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100110","11000101100001100101","11000101100001100101","11000101100001100101","11000101100001100101","11000101100001100101","11000101100001100101","11000101100001100101","11000101100001100101","11000101100001100101","11000101100001100101","11000101010001100101","11000101010001100101","11000101010001100101","11000101010001100101","11000101010001100101","11000101010001100101","11000101010001100101","11000101010001100101","11000101010001100101","11000101010001100101","11000101010001100101","11000101010001100101","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100100","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101010001100011","11000101000001100011","11000101000001100011","11000101000001100011","11000101000001100011","11000101000001100011","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100010","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100001","11000101000001100000","11000101000001100000","11000101000001100000","11000101000001100000","11000101000001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001100000","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011111","11000100110001011110","11000100110001011110","11000100110001011110","11000100110001011110","11000100110001011110","11000100110001011110","11000100110001011110","11000100110001011110","11000100110001011110","11000100110001011110","11000100110001011110","11000100110001011110","11000100110001011110","11000100110001011110","11000100110001011110","11000100100001011110","11000100100001011110","11000100100001011110","11000100100001011110","11000100100001011110","11000100100001011110","11000100100001011110","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011101","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011100","11000100100001011011","11000100100001011011","11000100100001011011","11000100100001011011","11000100100001011011","11000100100001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011011","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011010","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100010001011001","11000100000001011001","11000100000001011001","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001011000","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010111","11000100000001010110","11000100000001010110","11000100000001010110","11000100000001010110","11000100000001010110","11000100000001010110","11000100000001010110","11000100000001010110","11000100000001010110","11000100000001010110","11000100000001010110","11000100000001010110","11000100000001010110","11000100000001010110","11000011110001010110","11000011110001010110","11000011110001010110","11000011110001010110","11000011110001010110","11000011110001010110","11000011110001010110","11000011110001010110","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010101","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010100","11000011110001010011","11000011110001010011","11000011110001010011","11000011110001010011","11000011110001010011","11000011110001010011","11000011110001010011","11000011110001010011","11000011110001010011","11000011110001010011","11000011110001010011","11000011100001010011","11000011100001010011","11000011100001010011","11000011100001010011","11000011100001010011","11000011100001010011","11000011100001010011","11000011100001010011","11000011100001010011","11000011100001010011","11000011100001010011","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010010","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010001","11000011100001010000","11000011100001010000","11000011100001010000","11000011100001010000","11000011100001010000","11000011100001010000","11000011100001010000","11000011100001010000","11000011100001010000","11000011010001010000","11000011010001010000","11000011010001010000","11000011010001010000","11000011010001010000","11000011010001010000","11000011010001010000","11000011010001010000","11000011010001010000","11000011010001010000","11000011010001010000","11000011010001010000","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001111","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001110","11000011010001001101","11000011010001001101","11000011010001001101","11000011010001001101","11000011010001001101","11000011010001001101","11000011010001001101","11000011010001001101","11000011010001001101","11000011010001001101","11000011010001001101","11000011000001001101","11000011000001001101","11000011000001001101","11000011000001001101","11000011000001001101","11000011000001001101","11000011000001001101","11000011000001001101","11000011000001001101","11000011000001001101","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001100","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001011","11000011000001001010","11000011000001001010","11000011000001001010","11000011000001001010","11000011000001001010","11000011000001001010","11000011000001001010","11000011000001001010","11000011000001001010","11000011000001001010","11000011000001001010","11000011000001001010","11000011000001001010","11000011000001001010","11000011000001001010","11000011000001001010","11000010110001001010","11000010110001001010","11000010110001001010","11000010110001001010","11000010110001001010","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001001","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001001000","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000111","11000010110001000110","11000010110001000110","11000010110001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000110","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000101","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000100","11000010100001000011","11000010100001000011","11000010100001000011","11000010100001000011","11000010100001000011","11000010100001000011","11000010100001000011","11000010100001000011","11000010100001000011","11000010100001000011","11000010100001000011","11000010100001000011","11000010100001000011","11000010100001000011","11000010100001000011","11000010100001000011","11000010010001000011","11000010010001000011","11000010010001000011","11000010010001000011","11000010010001000011","11000010010001000011","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000010","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000001","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010001000000","11000010010000111111","11000010010000111111","11000010010000111111","11000010010000111111","11000010010000111111","11000010010000111111","11000010010000111111","11000010010000111111","11000010010000111111","11000010010000111111","11000010000000111111","11000010000000111111","11000010000000111111","11000010000000111111","11000010000000111111","11000010000000111111","11000010000000111111","11000010000000111111","11000010000000111111","11000010000000111111","11000010000000111111","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111110","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111101","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111100","11000010000000111011","11000010000000111011","11000010000000111011","11000010000000111011","11000010000000111011","11000010000000111011","11000010000000111011","11000010000000111011","11000010000000111011","11000010000000111011","11000010000000111011","11000001110000111011","11000001110000111011","11000001110000111011","11000001110000111011","11000001110000111011","11000001110000111011","11000001110000111011","11000001110000111011","11000001110000111011","11000001110000111011","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111010","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111001","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000111000","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001110000110111","11000001100000110111","11000001100000110111","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110110","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110101","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110100","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110011","11000001100000110010","11000001100000110010","11000001100000110010","11000001100000110010","11000001100000110010","11000001100000110010","11000001100000110010","11000001100000110010","11000001100000110010","11000001100000110010","11000001100000110010","11000001100000110010","11000001100000110010","11000001010000110010","11000001010000110010","11000001010000110010","11000001010000110010","11000001010000110010","11000001010000110010","11000001010000110010","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110001","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000110000","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101111","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101110","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001010000101101","11000001000000101101","11000001000000101101","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101100","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101011","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101010","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101001","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000101000","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000001000000100111","11000000110000100111","11000000110000100111","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100110","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100101","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100100","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100011","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100010","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100001","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000100000","11000000110000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011111","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011110","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011101","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011100","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011011","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011010","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011001","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000011000","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010111","11000000100000010110","11000000100000010110","11000000100000010110","11000000100000010110","11000000100000010110","11000000100000010110","11000000100000010110","11000000100000010110","11000000010000010110","11000000010000010110","11000000010000010110","11000000010000010110","11000000010000010110","11000000010000010110","11000000010000010110","11000000010000010110","11000000010000010110","11000000010000010110","11000000010000010110","11000000010000010110","11000000010000010110","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010101","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010100","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010011","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010010","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010001","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000010000","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001111","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001110","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001101","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001100","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001011","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001010","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001001","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000001000","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000111","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000110","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000101","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000100","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000011","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000010","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000001","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000000000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000010000000000","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111111","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111110","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111101","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111100","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111011","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111010","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111001","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111111000","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110111","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110110","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110101","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110100","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110011","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110010","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110001","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111110000","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101111","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101110","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101101","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101100","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101011","11000000011111101010","11000000011111101010","11000000011111101010","11000000011111101010","11000000011111101010","11000000011111101010","11000000011111101010","11000000011111101010","11000000011111101010","11000000011111101010","11000000011111101010","11000000011111101010","11000000011111101010","11000000101111101010","11000000101111101010","11000000101111101010","11000000101111101010","11000000101111101010","11000000101111101010","11000000101111101010","11000000101111101010","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101001","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111101000","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100111","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100110","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100101","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100100","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100011","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100010","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000101111100001","11000000111111100001","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111100000","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011111","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011110","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011101","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011100","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011011","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011010","11000000111111011001","11000000111111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011001","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111011000","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010111","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010110","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010101","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010100","11000001001111010011","11000001001111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010011","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010010","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010001","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111010000","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001111","11000001011111001110","11000001011111001110","11000001011111001110","11000001011111001110","11000001011111001110","11000001011111001110","11000001011111001110","11000001101111001110","11000001101111001110","11000001101111001110","11000001101111001110","11000001101111001110","11000001101111001110","11000001101111001110","11000001101111001110","11000001101111001110","11000001101111001110","11000001101111001110","11000001101111001110","11000001101111001110","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001101","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001100","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001011","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001010","11000001101111001001","11000001101111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001001","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111001000","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000111","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000110","11000001111111000101","11000001111111000101","11000001111111000101","11000001111111000101","11000001111111000101","11000001111111000101","11000001111111000101","11000001111111000101","11000001111111000101","11000001111111000101","11000010001111000101","11000010001111000101","11000010001111000101","11000010001111000101","11000010001111000101","11000010001111000101","11000010001111000101","11000010001111000101","11000010001111000101","11000010001111000101","11000010001111000101","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000100","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000011","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000010","11000010001111000001","11000010001111000001","11000010001111000001","11000010001111000001","11000010001111000001","11000010001111000001","11000010001111000001","11000010001111000001","11000010001111000001","11000010001111000001","11000010001111000001","11000010011111000001","11000010011111000001","11000010011111000001","11000010011111000001","11000010011111000001","11000010011111000001","11000010011111000001","11000010011111000001","11000010011111000001","11000010011111000001","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011111000000","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111111","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111110","11000010011110111101","11000010011110111101","11000010011110111101","11000010011110111101","11000010011110111101","11000010011110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111101","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111100","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111011","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010101110111010","11000010111110111010","11000010111110111010","11000010111110111010","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111001","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110111000","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110111","11000010111110110110","11000010111110110110","11000010111110110110","11000010111110110110","11000010111110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110110","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110101","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110100","11000011001110110011","11000011001110110011","11000011001110110011","11000011001110110011","11000011001110110011","11000011001110110011","11000011001110110011","11000011001110110011","11000011001110110011","11000011001110110011","11000011011110110011","11000011011110110011","11000011011110110011","11000011011110110011","11000011011110110011","11000011011110110011","11000011011110110011","11000011011110110011","11000011011110110011","11000011011110110011","11000011011110110011","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110010","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110001","11000011011110110000","11000011011110110000","11000011011110110000","11000011011110110000","11000011011110110000","11000011011110110000","11000011011110110000","11000011011110110000","11000011011110110000","11000011011110110000","11000011011110110000","11000011011110110000","11000011101110110000","11000011101110110000","11000011101110110000","11000011101110110000","11000011101110110000","11000011101110110000","11000011101110110000","11000011101110110000","11000011101110110000","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101111","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101110","11000011101110101101","11000011101110101101","11000011101110101101","11000011101110101101","11000011101110101101","11000011101110101101","11000011101110101101","11000011101110101101","11000011101110101101","11000011101110101101","11000011101110101101","11000011111110101101","11000011111110101101","11000011111110101101","11000011111110101101","11000011111110101101","11000011111110101101","11000011111110101101","11000011111110101101","11000011111110101101","11000011111110101101","11000011111110101101","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101100","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101011","11000011111110101010","11000011111110101010","11000011111110101010","11000011111110101010","11000011111110101010","11000011111110101010","11000011111110101010","11000011111110101010","11000100001110101010","11000100001110101010","11000100001110101010","11000100001110101010","11000100001110101010","11000100001110101010","11000100001110101010","11000100001110101010","11000100001110101010","11000100001110101010","11000100001110101010","11000100001110101010","11000100001110101010","11000100001110101010","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101001","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110101000","11000100001110100111","11000100001110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100111","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100110","11000100011110100101","11000100011110100101","11000100011110100101","11000100011110100101","11000100011110100101","11000100011110100101","11000100011110100101","11000100011110100101","11000100011110100101","11000100011110100101","11000100011110100101","11000100011110100101","11000100011110100101","11000100011110100101","11000100011110100101","11000100011110100101","11000100101110100101","11000100101110100101","11000100101110100101","11000100101110100101","11000100101110100101","11000100101110100101","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100100","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100011","11000100101110100010","11000100101110100010","11000100101110100010","11000100101110100010","11000100101110100010","11000100101110100010","11000100101110100010","11000100111110100010","11000100111110100010","11000100111110100010","11000100111110100010","11000100111110100010","11000100111110100010","11000100111110100010","11000100111110100010","11000100111110100010","11000100111110100010","11000100111110100010","11000100111110100010","11000100111110100010","11000100111110100010","11000100111110100010","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100001","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000100111110100000","11000101001110100000","11000101001110100000","11000101001110100000","11000101001110100000","11000101001110100000","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011111","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011110","11000101001110011101","11000101001110011101","11000101001110011101","11000101001110011101","11000101001110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011101","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011100","11000101011110011011","11000101011110011011","11000101011110011011","11000101011110011011","11000101011110011011","11000101011110011011","11000101011110011011","11000101011110011011","11000101011110011011","11000101011110011011","11000101011110011011","11000101011110011011","11000101101110011011","11000101101110011011","11000101101110011011","11000101101110011011","11000101101110011011","11000101101110011011","11000101101110011011","11000101101110011011","11000101101110011011","11000101101110011011","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011010","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101101110011001","11000101111110011001","11000101111110011001","11000101111110011001","11000101111110011001","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110011000","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010111","11000101111110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010110","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010101","11000110001110010100","11000110001110010100","11000110001110010100","11000110001110010100","11000110001110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010100","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010011","11000110011110010010","11000110011110010010","11000110011110010010","11000110011110010010","11000110011110010010","11000110011110010010","11000110011110010010","11000110101110010010","11000110101110010010","11000110101110010010","11000110101110010010","11000110101110010010","11000110101110010010","11000110101110010010","11000110101110010010","11000110101110010010","11000110101110010010","11000110101110010010","11000110101110010010","11000110101110010010","11000110101110010010","11000110101110010010","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010001","11000110101110010000","11000110101110010000","11000110101110010000","11000110101110010000","11000110101110010000","11000110101110010000","11000110101110010000","11000110101110010000","11000110101110010000","11000110111110010000","11000110111110010000","11000110111110010000","11000110111110010000","11000110111110010000","11000110111110010000","11000110111110010000","11000110111110010000","11000110111110010000","11000110111110010000","11000110111110010000","11000110111110010000","11000110111110010000","11000110111110010000","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001111","11000110111110001110","11000110111110001110","11000110111110001110","11000110111110001110","11000110111110001110","11000110111110001110","11000110111110001110","11000110111110001110","11000110111110001110","11000110111110001110","11000111001110001110","11000111001110001110","11000111001110001110","11000111001110001110","11000111001110001110","11000111001110001110","11000111001110001110","11000111001110001110","11000111001110001110","11000111001110001110","11000111001110001110","11000111001110001110","11000111001110001110","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001101","11000111001110001100","11000111001110001100","11000111001110001100","11000111001110001100","11000111001110001100","11000111001110001100","11000111001110001100","11000111001110001100","11000111001110001100","11000111011110001100","11000111011110001100","11000111011110001100","11000111011110001100","11000111011110001100","11000111011110001100","11000111011110001100","11000111011110001100","11000111011110001100","11000111011110001100","11000111011110001100","11000111011110001100","11000111011110001100","11000111011110001100","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001011","11000111011110001010","11000111011110001010","11000111011110001010","11000111011110001010","11000111011110001010","11000111011110001010","11000111011110001010","11000111011110001010","11000111101110001010","11000111101110001010","11000111101110001010","11000111101110001010","11000111101110001010","11000111101110001010","11000111101110001010","11000111101110001010","11000111101110001010","11000111101110001010","11000111101110001010","11000111101110001010","11000111101110001010","11000111101110001010","11000111101110001010","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001001","11000111101110001000","11000111101110001000","11000111101110001000","11000111101110001000","11000111101110001000","11000111101110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110001000","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000111","11000111111110000110","11000111111110000110","11000111111110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000110","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000001110000101","11001000011110000101","11001000011110000101","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000100","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000011110000011","11001000101110000011","11001000101110000011","11001000101110000011","11001000101110000011","11001000101110000011","11001000101110000011","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000010","11001000101110000001","11001000101110000001","11001000101110000001","11001000101110000001","11001000101110000001","11001000101110000001","11001000101110000001","11001000101110000001","11001000101110000001","11001000101110000001","11001000101110000001","11001000111110000001","11001000111110000001","11001000111110000001","11001000111110000001","11001000111110000001","11001000111110000001","11001000111110000001","11001000111110000001","11001000111110000001","11001000111110000001","11001000111110000001","11001000111110000001","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111110000000","11001000111101111111","11001000111101111111","11001000111101111111","11001000111101111111","11001000111101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111111","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001001101111110","11001001011101111110","11001001011101111110","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111101","11001001011101111100","11001001011101111100","11001001011101111100","11001001011101111100","11001001011101111100","11001001011101111100","11001001011101111100","11001001011101111100","11001001011101111100","11001001011101111100","11001001011101111100","11001001011101111100","11001001011101111100","11001001101101111100","11001001101101111100","11001001101101111100","11001001101101111100","11001001101101111100","11001001101101111100","11001001101101111100","11001001101101111100","11001001101101111100","11001001101101111100","11001001101101111100","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111011","11001001101101111010","11001001101101111010","11001001101101111010","11001001101101111010","11001001101101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111010","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001001111101111001","11001010001101111001","11001010001101111001","11001010001101111001","11001010001101111001","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101111000","11001010001101110111","11001010001101110111","11001010001101110111","11001010001101110111","11001010001101110111","11001010001101110111","11001010001101110111","11001010001101110111","11001010001101110111","11001010001101110111","11001010011101110111","11001010011101110111","11001010011101110111","11001010011101110111","11001010011101110111","11001010011101110111","11001010011101110111","11001010011101110111","11001010011101110111","11001010011101110111","11001010011101110111","11001010011101110111","11001010011101110111","11001010011101110111","11001010011101110111","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010011101110110","11001010101101110110","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110101","11001010101101110100","11001010101101110100","11001010101101110100","11001010101101110100","11001010101101110100","11001010101101110100","11001010101101110100","11001010101101110100","11001010101101110100","11001010101101110100","11001010101101110100","11001010101101110100","11001010111101110100","11001010111101110100","11001010111101110100","11001010111101110100","11001010111101110100","11001010111101110100","11001010111101110100","11001010111101110100","11001010111101110100","11001010111101110100","11001010111101110100","11001010111101110100","11001010111101110100","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001010111101110011","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110010","11001011001101110001","11001011001101110001","11001011001101110001","11001011001101110001","11001011001101110001","11001011001101110001","11001011001101110001","11001011001101110001","11001011001101110001","11001011001101110001","11001011001101110001","11001011001101110001","11001011001101110001","11001011011101110001","11001011011101110001","11001011011101110001","11001011011101110001","11001011011101110001","11001011011101110001","11001011011101110001","11001011011101110001","11001011011101110001","11001011011101110001","11001011011101110001","11001011011101110001","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011011101110000","11001011101101110000","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101111","11001011101101101110","11001011101101101110","11001011101101101110","11001011101101101110","11001011101101101110","11001011101101101110","11001011101101101110","11001011101101101110","11001011101101101110","11001011101101101110","11001011111101101110","11001011111101101110","11001011111101101110","11001011111101101110","11001011111101101110","11001011111101101110","11001011111101101110","11001011111101101110","11001011111101101110","11001011111101101110","11001011111101101110","11001011111101101110","11001011111101101110","11001011111101101110","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001011111101101101","11001100001101101101","11001100001101101101","11001100001101101101","11001100001101101101","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101100","11001100001101101011","11001100001101101011","11001100001101101011","11001100001101101011","11001100001101101011","11001100001101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101011","11001100011101101010","11001100011101101010","11001100011101101010","11001100011101101010","11001100011101101010","11001100011101101010","11001100011101101010","11001100011101101010","11001100011101101010","11001100011101101010","11001100011101101010","11001100011101101010","11001100011101101010","11001100011101101010","11001100011101101010","11001100011101101010","11001100101101101010","11001100101101101010","11001100101101101010","11001100101101101010","11001100101101101010","11001100101101101010","11001100101101101010","11001100101101101010","11001100101101101010","11001100101101101010","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100101101101001","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101101000","11001100111101100111","11001100111101100111","11001100111101100111","11001100111101100111","11001100111101100111","11001100111101100111","11001100111101100111","11001100111101100111","11001100111101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100111","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101001101100110","11001101011101100110","11001101011101100110","11001101011101100110","11001101011101100110","11001101011101100110","11001101011101100110","11001101011101100110","11001101011101100110","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101011101100101","11001101101101100101","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100100","11001101101101100011","11001101101101100011","11001101101101100011","11001101101101100011","11001101101101100011","11001101101101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100011","11001101111101100010","11001101111101100010","11001101111101100010","11001101111101100010","11001101111101100010","11001101111101100010","11001101111101100010","11001101111101100010","11001101111101100010","11001101111101100010","11001101111101100010","11001101111101100010","11001101111101100010","11001101111101100010","11001110001101100010","11001110001101100010","11001110001101100010","11001110001101100010","11001110001101100010","11001110001101100010","11001110001101100010","11001110001101100010","11001110001101100010","11001110001101100010","11001110001101100010","11001110001101100010","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110001101100001","11001110011101100001","11001110011101100001","11001110011101100001","11001110011101100001","11001110011101100001","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101100000","11001110011101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011111","11001110101101011110","11001110101101011110","11001110101101011110","11001110101101011110","11001110101101011110","11001110101101011110","11001110101101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011110","11001110111101011101","11001110111101011101","11001110111101011101","11001110111101011101","11001110111101011101","11001110111101011101","11001110111101011101","11001110111101011101","11001110111101011101","11001110111101011101","11001110111101011101","11001110111101011101","11001110111101011101","11001111001101011101","11001111001101011101","11001111001101011101","11001111001101011101","11001111001101011101","11001111001101011101","11001111001101011101","11001111001101011101","11001111001101011101","11001111001101011101","11001111001101011101","11001111001101011101","11001111001101011101","11001111001101011101","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111001101011100","11001111011101011100","11001111011101011100","11001111011101011100","11001111011101011100","11001111011101011100","11001111011101011100","11001111011101011100","11001111011101011100","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111011101011011","11001111101101011011","11001111101101011011","11001111101101011011","11001111101101011011","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011010","11001111101101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011001","11001111111101011000","11001111111101011000","11001111111101011000","11001111111101011000","11001111111101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101011000","11010000001101010111","11010000001101010111","11010000001101010111","11010000001101010111","11010000001101010111","11010000001101010111","11010000001101010111","11010000001101010111","11010000001101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010111","11010000011101010110","11010000011101010110","11010000011101010110","11010000011101010110","11010000011101010110","11010000011101010110","11010000011101010110","11010000011101010110","11010000011101010110","11010000011101010110","11010000011101010110","11010000011101010110","11010000101101010110","11010000101101010110","11010000101101010110","11010000101101010110","11010000101101010110","11010000101101010110","11010000101101010110","11010000101101010110","11010000101101010110","11010000101101010110","11010000101101010110","11010000101101010110","11010000101101010110","11010000101101010110","11010000101101010110","11010000101101010101","11010000101101010101","11010000101101010101","11010000101101010101","11010000101101010101","11010000101101010101","11010000101101010101","11010000101101010101","11010000101101010101","11010000101101010101","11010000101101010101","11010000101101010101","11010000101101010101","11010000101101010101","11010000101101010101","11010000101101010101","11010000111101010101","11010000111101010101","11010000111101010101","11010000111101010101","11010000111101010101","11010000111101010101","11010000111101010101","11010000111101010101","11010000111101010101","11010000111101010101","11010000111101010101","11010000111101010101","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010000111101010100","11010001001101010100","11010001001101010100","11010001001101010100","11010001001101010100","11010001001101010100","11010001001101010100","11010001001101010100","11010001001101010100","11010001001101010100","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001001101010011","11010001011101010011","11010001011101010011","11010001011101010011","11010001011101010011","11010001011101010011","11010001011101010011","11010001011101010011","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001011101010010","11010001101101010010","11010001101101010010","11010001101101010010","11010001101101010010","11010001101101010010","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001101101010001","11010001111101010001","11010001111101010001","11010001111101010001","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010001111101010000","11010010001101010000","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010001101001111","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010011101001110","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001101","11010010101101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001100","11010010111101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001011","11010011001101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011011101001010","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011101101001001","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010011111101001000","11010100001101001000","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100001101000111","11010100011101000111","11010100011101000111","11010100011101000111","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100011101000110","11010100101101000110","11010100101101000110","11010100101101000110","11010100101101000110","11010100101101000110","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100101101000101","11010100111101000101","11010100111101000101","11010100111101000101","11010100111101000101","11010100111101000101","11010100111101000101","11010100111101000101","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010100111101000100","11010101001101000100","11010101001101000100","11010101001101000100","11010101001101000100","11010101001101000100","11010101001101000100","11010101001101000100","11010101001101000100","11010101001101000100","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101001101000011","11010101011101000011","11010101011101000011","11010101011101000011","11010101011101000011","11010101011101000011","11010101011101000011","11010101011101000011","11010101011101000011","11010101011101000011","11010101011101000011","11010101011101000011","11010101011101000011","11010101011101000010","11010101011101000010","11010101011101000010","11010101011101000010","11010101011101000010","11010101011101000010","11010101011101000010","11010101011101000010","11010101011101000010","11010101011101000010","11010101011101000010","11010101011101000010","11010101011101000010","11010101011101000010","11010101011101000010","11010101011101000010","11010101101101000010","11010101101101000010","11010101101101000010","11010101101101000010","11010101101101000010","11010101101101000010","11010101101101000010","11010101101101000010","11010101101101000010","11010101101101000010","11010101101101000010","11010101101101000010","11010101101101000010","11010101101101000010","11010101101101000010","11010101101101000001","11010101101101000001","11010101101101000001","11010101101101000001","11010101101101000001","11010101101101000001","11010101101101000001","11010101101101000001","11010101101101000001","11010101101101000001","11010101101101000001","11010101101101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000001","11010101111101000000","11010101111101000000","11010101111101000000","11010101111101000000","11010101111101000000","11010101111101000000","11010101111101000000","11010101111101000000","11010101111101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001101000000","11010110001100111111","11010110001100111111","11010110001100111111","11010110001100111111","11010110001100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111111","11010110011100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110101100111110","11010110111100111110","11010110111100111110","11010110111100111110","11010110111100111110","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010110111100111101","11010111001100111101","11010111001100111101","11010111001100111101","11010111001100111101","11010111001100111101","11010111001100111101","11010111001100111101","11010111001100111101","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111001100111100","11010111011100111100","11010111011100111100","11010111011100111100","11010111011100111100","11010111011100111100","11010111011100111100","11010111011100111100","11010111011100111100","11010111011100111100","11010111011100111100","11010111011100111100","11010111011100111100","11010111011100111100","11010111011100111100","11010111011100111011","11010111011100111011","11010111011100111011","11010111011100111011","11010111011100111011","11010111011100111011","11010111011100111011","11010111011100111011","11010111011100111011","11010111011100111011","11010111011100111011","11010111011100111011","11010111011100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111011","11010111101100111010","11010111101100111010","11010111101100111010","11010111101100111010","11010111101100111010","11010111101100111010","11010111101100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111010","11010111111100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000001100111001","11011000011100111001","11011000011100111001","11011000011100111001","11011000011100111001","11011000011100111001","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000011100111000","11011000101100111000","11011000101100111000","11011000101100111000","11011000101100111000","11011000101100111000","11011000101100111000","11011000101100111000","11011000101100111000","11011000101100111000","11011000101100111000","11011000101100111000","11011000101100111000","11011000101100110111","11011000101100110111","11011000101100110111","11011000101100110111","11011000101100110111","11011000101100110111","11011000101100110111","11011000101100110111","11011000101100110111","11011000101100110111","11011000101100110111","11011000101100110111","11011000101100110111","11011000101100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110111","11011000111100110110","11011000111100110110","11011000111100110110","11011000111100110110","11011000111100110110","11011000111100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001001100110110","11011001011100110110","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001011100110101","11011001101100110101","11011001101100110101","11011001101100110101","11011001101100110101","11011001101100110101","11011001101100110101","11011001101100110101","11011001101100110101","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001101100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110100","11011001111100110011","11011001111100110011","11011001111100110011","11011001111100110011","11011001111100110011","11011001111100110011","11011001111100110011","11011001111100110011","11011001111100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010001100110011","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010011100110010","11011010101100110010","11011010101100110010","11011010101100110010","11011010101100110010","11011010101100110010","11011010101100110010","11011010101100110010","11011010101100110010","11011010101100110010","11011010101100110010","11011010101100110001","11011010101100110001","11011010101100110001","11011010101100110001","11011010101100110001","11011010101100110001","11011010101100110001","11011010101100110001","11011010101100110001","11011010101100110001","11011010101100110001","11011010101100110001","11011010101100110001","11011010101100110001","11011010101100110001","11011010101100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110001","11011010111100110000","11011010111100110000","11011010111100110000","11011010111100110000","11011010111100110000","11011010111100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011001100110000","11011011011100110000","11011011011100110000","11011011011100110000","11011011011100110000","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011011100101111","11011011101100101111","11011011101100101111","11011011101100101111","11011011101100101111","11011011101100101111","11011011101100101111","11011011101100101111","11011011101100101111","11011011101100101111","11011011101100101111","11011011101100101111","11011011101100101111","11011011101100101111","11011011101100101111","11011011101100101110","11011011101100101110","11011011101100101110","11011011101100101110","11011011101100101110","11011011101100101110","11011011101100101110","11011011101100101110","11011011101100101110","11011011101100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011011111100101110","11011100001100101110","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100001100101101","11011100011100101101","11011100011100101101","11011100011100101101","11011100011100101101","11011100011100101101","11011100011100101101","11011100011100101101","11011100011100101101","11011100011100101101","11011100011100101101","11011100011100101101","11011100011100101101","11011100011100101100","11011100011100101100","11011100011100101100","11011100011100101100","11011100011100101100","11011100011100101100","11011100011100101100","11011100011100101100","11011100011100101100","11011100011100101100","11011100011100101100","11011100011100101100","11011100011100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100101100101100","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011100111100101011","11011101001100101011","11011101001100101011","11011101001100101011","11011101001100101011","11011101001100101011","11011101001100101011","11011101001100101011","11011101001100101011","11011101001100101011","11011101001100101011","11011101001100101011","11011101001100101011","11011101001100101011","11011101001100101010","11011101001100101010","11011101001100101010","11011101001100101010","11011101001100101010","11011101001100101010","11011101001100101010","11011101001100101010","11011101001100101010","11011101001100101010","11011101001100101010","11011101001100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101011100101010","11011101101100101010","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101101100101001","11011101111100101001","11011101111100101001","11011101111100101001","11011101111100101001","11011101111100101001","11011101111100101001","11011101111100101001","11011101111100101001","11011101111100101001","11011101111100101001","11011101111100101001","11011101111100101001","11011101111100101001","11011101111100101001","11011101111100101001","11011101111100101000","11011101111100101000","11011101111100101000","11011101111100101000","11011101111100101000","11011101111100101000","11011101111100101000","11011101111100101000","11011101111100101000","11011101111100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110001100101000","11011110011100101000","11011110011100101000","11011110011100101000","11011110011100101000","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110011100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100111","11011110101100100110","11011110101100100110","11011110101100100110","11011110101100100110","11011110101100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011110111100100110","11011111001100100110","11011111001100100110","11011111001100100110","11011111001100100110","11011111001100100110","11011111001100100110","11011111001100100110","11011111001100100110","11011111001100100110","11011111001100100110","11011111001100100110","11011111001100100101","11011111001100100101","11011111001100100101","11011111001100100101","11011111001100100101","11011111001100100101","11011111001100100101","11011111001100100101","11011111001100100101","11011111001100100101","11011111001100100101","11011111001100100101","11011111001100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111011100100101","11011111101100100101","11011111101100100101","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111101100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100100","11011111111100100011","11011111111100100011","11011111111100100011","11011111111100100011","11011111111100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000001100100011","11100000011100100011","11100000011100100011","11100000011100100011","11100000011100100011","11100000011100100011","11100000011100100011","11100000011100100011","11100000011100100011","11100000011100100011","11100000011100100011","11100000011100100011","11100000011100100011","11100000011100100010","11100000011100100010","11100000011100100010","11100000011100100010","11100000011100100010","11100000011100100010","11100000011100100010","11100000011100100010","11100000011100100010","11100000011100100010","11100000011100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000101100100010","11100000111100100010","11100000111100100010","11100000111100100010","11100000111100100010","11100000111100100010","11100000111100100010","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100000111100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001001100100001","11100001011100100001","11100001011100100001","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001011100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100100000","11100001101100011111","11100001101100011111","11100001101100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100001111100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011111","11100010001100011110","11100010001100011110","11100010001100011110","11100010001100011110","11100010001100011110","11100010001100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010011100011110","11100010101100011110","11100010101100011110","11100010101100011110","11100010101100011110","11100010101100011110","11100010101100011110","11100010101100011110","11100010101100011110","11100010101100011110","11100010101100011110","11100010101100011110","11100010101100011110","11100010101100011110","11100010101100011110","11100010101100011110","11100010101100011101","11100010101100011101","11100010101100011101","11100010101100011101","11100010101100011101","11100010101100011101","11100010101100011101","11100010101100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100010111100011101","11100011001100011101","11100011001100011101","11100011001100011101","11100011001100011101","11100011001100011101","11100011001100011101","11100011001100011101","11100011001100011101","11100011001100011101","11100011001100011101","11100011001100011101","11100011001100011101","11100011001100011101","11100011001100011101","11100011001100011100","11100011001100011100","11100011001100011100","11100011001100011100","11100011001100011100","11100011001100011100","11100011001100011100","11100011001100011100","11100011001100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011011100011100","11100011101100011100","11100011101100011100","11100011101100011100","11100011101100011100","11100011101100011100","11100011101100011100","11100011101100011100","11100011101100011100","11100011101100011100","11100011101100011100","11100011101100011100","11100011101100011100","11100011101100011100","11100011101100011011","11100011101100011011","11100011101100011011","11100011101100011011","11100011101100011011","11100011101100011011","11100011101100011011","11100011101100011011","11100011101100011011","11100011101100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100011111100011011","11100100001100011011","11100100001100011011","11100100001100011011","11100100001100011011","11100100001100011011","11100100001100011011","11100100001100011011","11100100001100011011","11100100001100011011","11100100001100011011","11100100001100011011","11100100001100011011","11100100001100011011","11100100001100011011","11100100001100011010","11100100001100011010","11100100001100011010","11100100001100011010","11100100001100011010","11100100001100011010","11100100001100011010","11100100001100011010","11100100001100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100011100011010","11100100101100011010","11100100101100011010","11100100101100011010","11100100101100011010","11100100101100011010","11100100101100011010","11100100101100011010","11100100101100011010","11100100101100011010","11100100101100011010","11100100101100011010","11100100101100011010","11100100101100011010","11100100101100011010","11100100101100011010","11100100101100011001","11100100101100011001","11100100101100011001","11100100101100011001","11100100101100011001","11100100101100011001","11100100101100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100100111100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011001","11100101001100011000","11100101001100011000","11100101001100011000","11100101001100011000","11100101001100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101011100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100011000","11100101101100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100101111100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110001100010111","11100110011100010111","11100110011100010111","11100110011100010111","11100110011100010111","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110011100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110101100010110","11100110111100010110","11100110111100010110","11100110111100010110","11100110111100010110","11100110111100010110","11100110111100010110","11100110111100010110","11100110111100010110","11100110111100010110","11100110111100010110","11100110111100010101","11100110111100010101","11100110111100010101","11100110111100010101","11100110111100010101","11100110111100010101","11100110111100010101","11100110111100010101","11100110111100010101","11100110111100010101","11100110111100010101","11100110111100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111001100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010101","11100111011100010100","11100111011100010100","11100111011100010100","11100111011100010100","11100111011100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111101100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11100111111100010100","11101000001100010100","11101000001100010100","11101000001100010100","11101000001100010100","11101000001100010100","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000001100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000011100010011","11101000101100010011","11101000101100010011","11101000101100010011","11101000101100010011","11101000101100010011","11101000101100010011","11101000101100010011","11101000101100010011","11101000101100010011","11101000101100010011","11101000101100010011","11101000101100010011","11101000101100010011","11101000101100010011","11101000101100010011","11101000101100010010","11101000101100010010","11101000101100010010","11101000101100010010","11101000101100010010","11101000101100010010","11101000101100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101000111100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001001100010010","11101001011100010010","11101001011100010010","11101001011100010010","11101001011100010010","11101001011100010010","11101001011100010010","11101001011100010001","11101001011100010001","11101001011100010001","11101001011100010001","11101001011100010001","11101001011100010001","11101001011100010001","11101001011100010001","11101001011100010001","11101001011100010001","11101001011100010001","11101001011100010001","11101001011100010001","11101001011100010001","11101001011100010001","11101001011100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001101100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010001","11101001111100010000","11101001111100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010001100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010011100010000","11101010101100010000","11101010101100010000","11101010101100010000","11101010101100010000","11101010101100010000","11101010101100010000","11101010101100010000","11101010101100010000","11101010101100010000","11101010101100010000","11101010101100010000","11101010101100010000","11101010101100010000","11101010101100010000","11101010101100001111","11101010101100001111","11101010101100001111","11101010101100001111","11101010101100001111","11101010101100001111","11101010101100001111","11101010101100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101010111100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011001100001111","11101011011100001111","11101011011100001111","11101011011100001111","11101011011100001111","11101011011100001111","11101011011100001111","11101011011100001111","11101011011100001111","11101011011100001111","11101011011100001111","11101011011100001111","11101011011100001110","11101011011100001110","11101011011100001110","11101011011100001110","11101011011100001110","11101011011100001110","11101011011100001110","11101011011100001110","11101011011100001110","11101011011100001110","11101011011100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011101100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101011111100001110","11101100001100001110","11101100001100001110","11101100001100001110","11101100001100001110","11101100001100001110","11101100001100001110","11101100001100001110","11101100001100001110","11101100001100001110","11101100001100001101","11101100001100001101","11101100001100001101","11101100001100001101","11101100001100001101","11101100001100001101","11101100001100001101","11101100001100001101","11101100001100001101","11101100001100001101","11101100001100001101","11101100001100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100011100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100101100001101","11101100111100001101","11101100111100001101","11101100111100001101","11101100111100001101","11101100111100001101","11101100111100001101","11101100111100001101","11101100111100001101","11101100111100001101","11101100111100001101","11101100111100001101","11101100111100001100","11101100111100001100","11101100111100001100","11101100111100001100","11101100111100001100","11101100111100001100","11101100111100001100","11101100111100001100","11101100111100001100","11101100111100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101001100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101011100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001100","11101101101100001011","11101101101100001011","11101101101100001011","11101101101100001011","11101101101100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101101111100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110001100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110011100001011","11101110101100001011","11101110101100001011","11101110101100001011","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110101100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101110111100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111001100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001010","11101111011100001001","11101111011100001001","11101111011100001001","11101111011100001001","11101111011100001001","11101111011100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111101100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11101111111100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000001100001001","11110000011100001001","11110000011100001001","11110000011100001001","11110000011100001001","11110000011100001001","11110000011100001001","11110000011100001001","11110000011100001001","11110000011100001001","11110000011100001001","11110000011100001000","11110000011100001000","11110000011100001000","11110000011100001000","11110000011100001000","11110000011100001000","11110000011100001000","11110000011100001000","11110000011100001000","11110000011100001000","11110000011100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000101100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110000111100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001001100001000","11110001011100001000","11110001011100001000","11110001011100001000","11110001011100001000","11110001011100001000","11110001011100001000","11110001011100001000","11110001011100001000","11110001011100001000","11110001011100001000","11110001011100001000","11110001011100000111","11110001011100000111","11110001011100000111","11110001011100000111","11110001011100000111","11110001011100000111","11110001011100000111","11110001011100000111","11110001011100000111","11110001011100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001101100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110001111100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010001100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000111","11110010011100000110","11110010011100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010101100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110010111100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011001100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011011100000110","11110011101100000110","11110011101100000110","11110011101100000110","11110011101100000110","11110011101100000110","11110011101100000110","11110011101100000110","11110011101100000110","11110011101100000110","11110011101100000110","11110011101100000110","11110011101100000110","11110011101100000110","11110011101100000101","11110011101100000101","11110011101100000101","11110011101100000101","11110011101100000101","11110011101100000101","11110011101100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110011111100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100001100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100011100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100101100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000101","11110100111100000100","11110100111100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101001100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101011100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101101100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110101111100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110001100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000100","11110110011100000011","11110110011100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110101100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110110111100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111001100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111011100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111101100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11110111111100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000001100000011","11111000011100000011","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000011100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000101100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111000111100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001001100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001011100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001101100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111001111100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010001100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010011100000010","11111010101100000010","11111010101100000010","11111010101100000010","11111010101100000010","11111010101100000010","11111010101100000010","11111010101100000010","11111010101100000010","11111010101100000001","11111010101100000001","11111010101100000001","11111010101100000001","11111010101100000001","11111010101100000001","11111010101100000001","11111010101100000001","11111010101100000001","11111010101100000001","11111010101100000001","11111010101100000001","11111010101100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111010111100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011001100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011011100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011101100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111011111100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100001100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100011100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100101100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111100111100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101001100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101011100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101101100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111101111100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110001100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110011100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110101100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111110111100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111001100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111011100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111101100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","11111111111100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001","00000000001100000001");
begin
   process(clk)   begin       if (rising_edge(clk)) then           value <= rom_mem(to_integer(unsigned(addr)));
       end if;   end process;end rom_b;
