library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    generic(
        width :integer:=12;
        length :integer
    ) ;
    port (
        addr: in std_logic_vector(length-1 downto 0);
        value: out std_logic_vector(width-1 downto 0)
    );
end rom;

architecture rom_b of rom is
    type MEMORY is array(0 to 3) of std_logic_vector(width-1 downto 0);
    signal rom_mem :MEMORY :=(
        "000000010000","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111111001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111110001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111101001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111100001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001111","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111011001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111010001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001110","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111001001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","111000001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001101","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110111001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001100","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110110001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001011","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110101001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001010","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110100001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001001","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011001000","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110011000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000111","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000110","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110010000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000101","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000100","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000011","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000010","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000001","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110000000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001000000","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111111","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111110","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111101","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111100","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110001111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111011","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111010","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110010111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111001","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011111000","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110011110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110111","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110100110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110110","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110101110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110101","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110110110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110100","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","110111110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111000110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110011","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111001110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111010110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110010","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111011110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111100110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111101110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111110110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","111111110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110000","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000000110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000001110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000010110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000011110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000100110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110001","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000101110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000110110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110010","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","000111110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001000110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110011","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001001110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110100","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001010110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110101","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001011110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110110","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001100110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101110111","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111000","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001101111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111001","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111010","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001110111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111011","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111100","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111101","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111110","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111111111","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","010000000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000000","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000001","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000010","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000011","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000100","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001111000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000101","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000110","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001110000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101000111","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001000","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001101001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001001","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001100001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001010","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001011001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001011","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001010001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001100","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001001001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","001000001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001101","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000111001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000110001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001110","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000101001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000100001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000011001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000010001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000001001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111","000000001111"
);
begin


    value <= rom_mem(to_integer(unsigned(addr)));

end rom_b;