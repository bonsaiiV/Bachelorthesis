library ieee;
use ieee.std_logic_1164.all;
entity fft_tb is
end fft_tb;
architecture test of fft_tb is
    component fft
    generic(N : integer;
            width :integer; 
            width_twiddle : integer);
    port (
       clk, fft_start: in std_logic;
       output_valid : out std_logic;
       inA, inB : std_logic_vector(2*width-1 downto 0);
       outA, outB: std_logic_vector(2*width-1 downto 0));
    end component;
    signal clk, fft_start : std_logic := '0';
    signal inA, inB : std_logic_vector(37 downto 0) := (others =>'0');
    signal output_valid : std_logic;
    signal outA, outB : std_logic_vector(37 downto 0);
begin
    fft_i: fft
    generic map (
        width => 19,
        width_twiddle => 6,
        N => 15
    )
    port map (
        clk => clk,
        fft_start => fft_start,
        inA => inA,
        inB => inB,
        fft_done => fft_done,
        outA => outA,
        outB => outB
    );
   process begin
        wait for 1 ns;
        clk <= '1';
        wait for 1 ns;
        clk <= '0';
        fft_start <= '1';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000100100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110001110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000100010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000000111110101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101111110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000000111110101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000100101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000100011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000101100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000110000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111110100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101111010000000";
inB<="00000000000000000001000100000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000100110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000011111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111110010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111110100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100011010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000100000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111110100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000000111110111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000000111110111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100101110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111110011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000100011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100110010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111110111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101001000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111110111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000100001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000000111110111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100111010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111110100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000100011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111101100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000011111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101000010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000011111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111110010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110000100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000100100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000011111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110000000000";
inB<="00000000000000000001000100111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111110100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000000111110101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111110001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000100001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110000000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111110101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111101110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111110111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000100110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100101000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000000111101111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000100010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000101010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000100011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000011111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000100001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111110101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111110010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000100010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111110111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111110000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110000000000";
inB<="00000000000000000000111110010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000000111110100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000100111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000100001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111110010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010110000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000000111110001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111100000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000100101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000100001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101001100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000100011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000011110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110001110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111101110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101011100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110000100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000100001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000011111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110000110000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000100010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000100101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111110000000";
inB<="00000000000000000001000011111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111110101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100111100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111110110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111110110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111110110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111110101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110001100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000101000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000011110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101110010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000100011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000100101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000100110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111110100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100100000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000100010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101001110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111110010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111110010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111110111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000100000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000100010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000011111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100101100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100111000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000011110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000100010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000100010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000011110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011100000000";
inB<="00000000000000000001000100011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111110100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101001010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000100111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111110100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000100100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100011110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000100101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111110101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101010000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111110100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001000000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000100001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000000111110111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000101010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111110101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101101000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111110011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000100010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000100100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000100110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000011110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111110001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101111110000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000100001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000100010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000000111110011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100011110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111110100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110001000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000100011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000000111110101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000000111110111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100111010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000100001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110001100000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110000000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000100000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111110011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000000111110100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011010000000";
inB<="00000000000000000001000100011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000000111110111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000100010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000100000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000100001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000011110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000100100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000100001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000000111110110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111110001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111101110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111110111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000100110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000100010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000011111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110000000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111110110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111110001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100101000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111110011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000011111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000101011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111110100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000100011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000011111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000100010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111100000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111110101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101000010000000";
inB<="00000000000000000000111110001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101011010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111110001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100101100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100101010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101011110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100101100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000000111110101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111110010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000011111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110000110000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111110111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000100101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000100110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111110011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010010000000";
inB<="00000000000000000000111110010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000100001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111110111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101010100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111110101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111110100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011010000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111110100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000011111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000100000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000000111110110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101000100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000100101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110001100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000100001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000100010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000000111110001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000100110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111101011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111110101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010000000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111110100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000110010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000100011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111110111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000100100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111110101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111110010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000100001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100101110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101001010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111110111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000101011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000100001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101110010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000100011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100011010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111110010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000011111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000011111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010000000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100011010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000100010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100101010000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000100110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110001010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000011111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000000111110011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111110100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111110111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000100010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111110101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000101000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101000100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101010000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101100100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000100110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111101111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111110000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000100011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111110100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101111110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000100111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000100011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110001110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110001000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000100000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111101000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000100000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111110000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101101000000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000000111110100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111110100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111110000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100111000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000000111110111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101010010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100011010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000000111110101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000100101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111110101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101110110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100011010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101010000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000100001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111101111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000100110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100011010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000100000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110000010000000";
inB<="00000000000000000001000101101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000100000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101111000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111100110110000000";
inB<="00000000000000000001000100001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101101010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111110111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111110111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000000111101111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000011110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111110000000";
inB<="00000000000000000000111101111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100110010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100110000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011100000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000100001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111110111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000100010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000000111110101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000100110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000100101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111110100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111100000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000100001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000100000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111110111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100011110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000100011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100011110000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100111000000000";
inB<="00000000000000000000111110111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111110111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000000111110100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100000000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111101110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111110111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000100010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101001000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110001000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101011000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111110110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111101000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111010000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110000010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000100010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000011111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000000111110010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000100001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100110010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100011000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111110011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000000111110101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000100101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000011111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111110111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100101000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000100011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000100000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110010000000";
inB<="00000000000000000001000100100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101001000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000100110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000011110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101100100000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000100101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000000111110110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000101011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100110010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111110011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000100010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101110010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000000111110100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000100111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000100000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000000111110100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110001110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000000111110111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000000111110010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111110011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000000111110111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111110101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100101100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000100101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011110000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111110000000";
inB<="00000000000000000000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111110001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111110011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100111100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000100001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110001100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101111000000000";
inB<="00000000000000000000111110101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111110011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000100000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000100010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000100000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100011110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000000111110111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000100000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000100000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000100010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100110000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111110011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111110110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111110111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000101001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010110000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111110010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000100111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000100101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000000111110110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000100101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000100001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111110011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111110000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110001110000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110000000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100010000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000100001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000000111110100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111110001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000100010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000110000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000011111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000100011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111110011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111101111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111000000000";
inB<="00000000000000000001000100101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001010000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000000111110110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000000111101111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100000000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101100010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111110011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000100000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000100000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110010000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111110111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111110110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101010010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000000111101110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000011111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111100110000000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000100110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101101010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110100110000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000100011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000100000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111101101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000100010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100101110000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000011101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111110010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101000000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000000111110111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000100001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101011010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000011100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000100101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100110110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000101000000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111100000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100010000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111000110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000100100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000100010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111110110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000100011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000110000000";
inB<="00000000000000000000111111001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101110100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111010000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000011111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000011010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000000111111000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111110011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100010000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000011011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000100011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000100001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000011110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000100000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000100000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101010000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000000111110111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100001100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000100101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000011000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011111000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000000111110101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110010000000";
inB<="00000000000000000001000011110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111110110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000011100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000011000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010000000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110110000000";
inB<="00000000000000000000111111100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000000111111001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000100000000";
inB<="00000000000000000001000011001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000000111111001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001010000000";
inB<="00000000000000000001000101000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110111010000000";
inB<="00000000000000000000111111110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011000000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010000000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000011100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000010000000";
inB<="00000000000000000001000010101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010100000000";
inB<="00000000000000000001000010100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000100110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000001010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000011101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111100000000";
inB<="00000000000000000001000011111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000000111110111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001100000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000000111110010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000100000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111101101000000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011010000000";
inB<="00000000000000000000111111000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000011010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000011010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000011110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110100000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000011011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101010000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011010000000";
inB<="00000000000000000000111110100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001110000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000000111110110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100000000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000000111111010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000010111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111110000000";
inB<="00000000000000000001000011010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111110111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010110000000";
inB<="00000000000000000001000010111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110110110000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010010000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110110000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001010000000";
inB<="00000000000000000001000000101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110110000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000100000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000000111110111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000100001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110000000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000000111111010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000000110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000001000011001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000001000000111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000000111111101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011001000000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000011101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110010110000000";
inB<="00000000000000000001000001010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000000100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000000100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111100000000";
inB<="00000000000000000001000011001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110101100000000";
inB<="00000000000000000001000001111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111000000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100010000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000110000000";
inB<="00000000000000000001000010100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000001110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100000000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111111010000000";
inB<="00000000000000000001000011000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000000111111100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000110000000";
inB<="00000000000000000001000001101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011110000000";
inB<="00000000000000000001000000111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001010000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100110000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000010010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100100100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011110010000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110010000000";
inB<="00000000000000000001000001101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000100000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000000111111111010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000010101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010100000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000000000000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011000000000";
inB<="00000000000000000001000001000010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000010000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101000000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000000000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110100000000";
inB<="00000000000000000001000010110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101100000000";
inB<="00000000000000000001000010101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000001001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000000111111111110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010000000000";
inB<="00000000000000000001000010110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111110011100000000";
inB<="00000000000000000001000011111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011100000000";
inB<="00000000000000000001000000001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011100110000000";
inB<="00000000000000000001000000001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000010000110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111100100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101110000000";
inB<="00000000000000000001000010011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000000000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111010000000";
inB<="00000000000000000001000011011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000001000001100110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011010110000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001000000000";
inB<="00000000000000000001000010011110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111110000000000";
inB<="00000000000000000001000000110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101000000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111110000000";
inB<="00000000000000000001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110100000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111011110000000";
inB<="00000000000000000000111111100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111010110000000";
inB<="00000000000000000001000100111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011110000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000000111111101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100010000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011000000000";
inB<="00000000000000000001000010011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000001000000011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010110000000";
inB<="00000000000000000001000010100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000010110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000110100000000";
inB<="00000000000000000001000001001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000100110000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000001111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001000000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010010000000";
inB<="00000000000000000001000001101110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110110000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111110000000";
inB<="00000000000000000001000001001110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011011100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000001000000011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001100000000";
inB<="00000000000000000001000001100010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111010000000";
inB<="00000000000000000001000000101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000000111111001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000000110100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101000000000";
inB<="00000000000000000001000010010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000000111111110110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000100000000000000";
inB<="00000000000000000000111111011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010110000000";
inB<="00000000000000000001000010001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001010000000";
inB<="00000000000000000001000001010100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000011100000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000010011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000011101000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111100000000";
inB<="00000000000000000001000001010000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111101110000000";
inB<="00000000000000000000111110111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010100110000000";
inB<="00000000000000000001000010001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000001110000000";
inB<="00000000000000000000111110010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101010000000";
inB<="00000000000000000001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101100000000";
inB<="00000000000000000001000001110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011100000000";
inB<="00000000000000000001000010001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101000000000";
inB<="00000000000000000000111111111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001110010000000";
inB<="00000000000000000001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001100110000000";
inB<="00000000000000000001000000101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010000000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000100000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010010100000000";
inB<="00000000000000000001000001100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010100000000";
inB<="00000000000000000000111111110000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010110000000000";
inB<="00000000000000000001000000010110000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001100000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000111000000000";
inB<="00000000000000000001000001011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000000111111001000000000";
inB<="00000000000000000001000010010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000010010000000";
inB<="00000000000000000001000001110010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001000000000";
inB<="00000000000000000001000000010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001101110000000";
inB<="00000000000000000001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001100000000";
inB<="00000000000000000000111111011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111110000000";
inB<="00000000000000000001000000100100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101010000000";
inB<="00000000000000000001000001011000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111110111000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011101110000000";
inB<="00000000000000000001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001011000000000";
inB<="00000000000000000000111111101100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010000000000000";
inB<="00000000000000000001000001000100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001000000000000";
inB<="00000000000000000000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010111010000000";
inB<="00000000000000000000111111111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010011110000000";
inB<="00000000000000000000111111010010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001010010000000";
inB<="00000000000000000001000000001100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000011000110000000";
inB<="00000000000000000001000000111100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010101100000000";
inB<="00000000000000000001000000001000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001111000000000";
inB<="00000000000000000001000000011100000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000010001010000000";
inB<="00000000000000000001000001011010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000000101110000000";
inB<="00000000000000000001000011001010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="00000000000000000001000001001110000000";
inB<="00000000000000000001000001101010000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
while output_valid = '0' loop
            wait for 1 ns;
            clk <= '1';
            wait for 1 ns;
            clk <= '0';
        end loop;
        for i in 0 to 16500 loop
        wait for 1 ns;
            clk <= '1';
            wait for 1 ns;
            clk <= '0';
        end loop;
        wait;
    end process;
end test;
