library ieee;
use ieee.std_logic_1164.all;
entity fft_tb is
end fft_tb;
architecture test of fft_tb is
    component fft
    port (
       clk, fft_start: in std_logic;
       output_valid : out std_logic;
       inA, inB : in std_logic_vector(47 downto 0);
       outA, outB: out std_logic_vector(47 downto 0));
    end component;
signal inA, inB, outA, outB : std_logic_vector(47 downto 0) := (others =>'0');
    signal clk, fft_start : std_logic := '0';
    signal output_valid : std_logic;
begin
    fft_i: fft
    port map (
        clk => clk,
        fft_start => fft_start,
        inA => inA,
        inB => inB,
        output_valid => output_valid,
        outA => outA,
        outB => outB
    );
   process begin
        wait for 1 ns;
        clk <= '1';
        wait for 1 ns;
        clk <= '0';
        fft_start <= '1';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010001001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100011100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100101100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000001111101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000010100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011111100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001000100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000001111101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010001001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010001000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010001011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100110000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011110100000000000";
inB<="000000000000000000000000010001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100111000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000110100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000001111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000001111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001011100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010001000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001100100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100110100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111010010000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100101000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000001111101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100101000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001110100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010001000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100100100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010000100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100001000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010001001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100000000000000";
inB<="000000000000000000000000010001001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000001111101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100111000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100000000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010001001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001010000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000001111011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010001010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010001000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100000000000000";
inB<="000000000000000000000000001111100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000001111101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010001001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000101100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000001111100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000101100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101001100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000101100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010001000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100011100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100110100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010111000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100101100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100001100000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001000000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101000100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010001001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111100000000000";
inB<="000000000000000000000000010000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001111000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100011000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010001010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011100100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010001001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010001001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000101000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101001000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010011100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010001000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001011000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001110000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100111000000000000";
inB<="000000000000000000000000010001000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010010100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010001001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010001001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100111000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001000000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000111100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010001001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000010000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000001111101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010001010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011010000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010001000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010001001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000010100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000010000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010001001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011111100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010001000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101000100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000001111100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000111100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100010000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010001000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000001111101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000101100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000001111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001110100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100011000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101001000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100000000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000001111101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100110100000000000";
inB<="000000000000000000000000010001000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000001111101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010001000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010001001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000001111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010001001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000010000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100000000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000101100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001010000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010001010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010001000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100111100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010000100000000000";
inB<="000000000000000000000000001111100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111010110100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001011000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001010100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010111100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001000000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001011000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000001111101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100001100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010001001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100110100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010001001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101000100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100100000000000";
inB<="000000000000000000000000001111100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111010101000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100110100000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000101100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101000000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100101000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000001111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010001000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010001001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100011000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000001111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010001001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000010100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010001100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010001000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101001000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010001001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000010000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001011100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111010010100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010001010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011100100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010001000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000110100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101001100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100100000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000110100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010001000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001010100000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010001001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000010100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100010100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000001111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010001000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010001010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010001000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010100000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011001000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010001001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010001000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100110000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011111100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010001001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010001000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100011100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100010000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101001000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011010000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000001111101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001110000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000001111101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111010100100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000110100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000001111101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011101100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000110100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000001111100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010100000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010001001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000110100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100101100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101001000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000001111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100000100000000000";
inB<="000000000000000000000000010001011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011110000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111001101100000000000";
inB<="000000000000000000000000010001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011010100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000001111011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111100000000000";
inB<="000000000000000000000000001111011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001100100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100111000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101001100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010001000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000001111101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010001001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010001001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000111100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000101000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010001000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000111100000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001110000000000000";
inB<="000000000000000000000000001111101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000001111101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001000000000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100010000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010110000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100000100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010001010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001000100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000001111100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010001000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100101000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001100100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000110000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000001111101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001000100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010001000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100111000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100110100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100100000000000";
inB<="000000000000000000000000010001001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010010000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010001001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011001000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010001001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000001111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100110100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010001010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001100100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100110000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011100100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000010000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000001111101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010001001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000001111101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100011100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000001111101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000001111100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000001111101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001011000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010001001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010001001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100111100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111100000000000";
inB<="000000000000000000000000001111101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001111000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001000000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011110000000000000";
inB<="000000000000000000000000001111101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010001000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000111100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000001111101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111111000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010001000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001100000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010001010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100101100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010001001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010001001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000001111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010001001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010001000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100011100000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000100000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010001000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000001111101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101010000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010001000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101000100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100111000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110000000000000";
inB<="000000000000000000000000010001001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000010100000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000001111101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000001111011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001000000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011000100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010001000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000001111011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111001100000000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010001001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100110100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001011010100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101001100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010001000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001000000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010001000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001011100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110000100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001000100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010000000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111101000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000001111101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111010110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010001001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001010000000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111000000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111000100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110001100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010001001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010001000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101111100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010001000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000001100000000000";
inB<="000000000000000000000000001111110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011101000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110100000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000001111110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000110111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010001000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010001000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010001000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000001111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000011000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010001001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000110001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111110000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000001111101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101100100000000000";
inB<="000000000000000000000000010000111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110110100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111111011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000110000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100000000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101100000000000";
inB<="000000000000000000000000001111111001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110000000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000001111110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001000000000000";
inB<="000000000000000000000000010000110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000001111110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010100000000000";
inB<="000000000000000000000000010001010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101110100000000000";
inB<="000000000000000000000000001111111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000010001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110110000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000100000000000";
inB<="000000000000000000000000010000101011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101000000000000";
inB<="000000000000000000000000010000101000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010001001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000010101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111000000000000";
inB<="000000000000000000000000010000111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000001111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110011000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000001111110000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000001111100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010001000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111011010000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000011111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110100000000000";
inB<="000000000000000000000000001111110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000110100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000111101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111000000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100111000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110100000000000";
inB<="000000000000000000000000001111101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000001111101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001000000000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000101010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000001111110101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111111100000000000";
inB<="000000000000000000000000010000110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111101111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101100000000000";
inB<="000000000000000000000000010000101110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101101100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110100100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101100000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000001110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010100000000000";
inB<="000000000000000000000000010000001010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101100000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001000000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000001111101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010001000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100000000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000001111110101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000001100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000101111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000010000110011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000000000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000010000001110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000001111111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110010000000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000111010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000011010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100101100000000000";
inB<="000000000000000000000000010000010100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000001001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000001000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000011101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111000000000000";
inB<="000000000000000000000000010000110011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111101011000000000000";
inB<="000000000000000000000000010000011111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000100000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110000000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000100000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000001100000000000";
inB<="000000000000000000000000010000101001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000011101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011000000000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111110100000000000";
inB<="000000000000000000000000010000110001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000001111111001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001100000000000";
inB<="000000000000000000000000010000011011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111100000000000";
inB<="000000000000000000000000010000001111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000100100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001001001000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110100100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111100100000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001100100000000000";
inB<="000000000000000000000000010000011010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010001000000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000001111111110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000101011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000000000000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000110000000000000";
inB<="000000000000000000000000010000010000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000100000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101010000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010000000001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111101000000000000";
inB<="000000000000000000000000010000101100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011000000000000";
inB<="000000000000000000000000010000101010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000010011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000001111111111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100000000000000";
inB<="000000000000000000000000010000101101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111100111000000000000";
inB<="000000000000000000000000010000111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111000000000000";
inB<="000000000000000000000000010000000011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111001100000000000";
inB<="000000000000000000000000010000000010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000100001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111001000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011100000000000";
inB<="000000000000000000000000010000100110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000000001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110100000000000";
inB<="000000000000000000000000010000110110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000010000011001100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110101100000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010000000000000";
inB<="000000000000000000000000010000100111100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111100000000000000";
inB<="000000000000000000000000010000001101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001010000000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111100000000000";
inB<="000000000000000000000000010000011000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101101000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110111100000000000";
inB<="000000000000000000000000001111111000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110101100000000000";
inB<="000000000000000000000000010001001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111100000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000001111111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101000100000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100110000000000000";
inB<="000000000000000000000000010000100111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000010000000110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000010000001000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101100000000000";
inB<="000000000000000000000000010000101001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000101100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001101000000000000";
inB<="000000000000000000000000010000010010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001001100000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000011110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010000000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100100100000000000";
inB<="000000000000000000000000010000011011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011101100000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011111100000000000";
inB<="000000000000000000000000010000010011100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000010000000110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110011000000000000";
inB<="000000000000000000000000010000011000100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000001100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110100000000000";
inB<="000000000000000000000000010000001010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000001111110010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000001101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111010000000000000";
inB<="000000000000000000000000010000100101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000001111111101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010001000000000000000000";
inB<="000000000000000000000000001111110110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010101100000000000";
inB<="000000000000000000000000010000100011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000010100000000000";
inB<="000000000000000000000000010000010101000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000111000000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000100110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000111010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001111000000000000";
inB<="000000000000000000000000010000010100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111111011100000000000";
inB<="000000000000000000000000001111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101001100000000000";
inB<="000000000000000000000000010000100010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000011100000000000";
inB<="000000000000000000000000001111100101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111111100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010100000000000";
inB<="000000000000000000000000010000010000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011000000000000";
inB<="000000000000000000000000010000011100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010111000000000000";
inB<="000000000000000000000000010000100010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011010000000000000";
inB<="000000000000000000000000001111111110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000010010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011100100000000000";
inB<="000000000000000000000000010000000000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011001100000000000";
inB<="000000000000000000000000010000001011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100000000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100001000000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100101000000000000";
inB<="000000000000000000000000010000011001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000101000000000000";
inB<="000000000000000000000000001111111100000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101100000000000000";
inB<="000000000000000000000000010000000101100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100011000000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001110000000000000";
inB<="000000000000000000000000010000010111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000001111110010000000000000";
inB<="000000000000000000000000010000100100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000000100100000000000";
inB<="000000000000000000000000010000011100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010010000000000000";
inB<="000000000000000000000000010000000100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011011100000000000";
inB<="000000000000000000000000010000101000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011000000000000";
inB<="000000000000000000000000001111110111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101111100000000000";
inB<="000000000000000000000000010000001001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111010100000000000";
inB<="000000000000000000000000010000010110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111101110000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000111011100000000000";
inB<="000000000000000000000000010000100000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010110000000000000";
inB<="000000000000000000000000001111111011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100000000000000000";
inB<="000000000000000000000000010000010001000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010000000000000000";
inB<="000000000000000000000000001111111000000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101110100000000000";
inB<="000000000000000000000000001111111111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100111100000000000";
inB<="000000000000000000000000001111110100100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010100100000000000";
inB<="000000000000000000000000010000000011000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000110001100000000000";
inB<="000000000000000000000000010000001111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000101011000000000000";
inB<="000000000000000000000000010000000010000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000011110000000000000";
inB<="000000000000000000000000010000000111000000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000100010100000000000";
inB<="000000000000000000000000010000010110100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000001011100000000000";
inB<="000000000000000000000000010000110010100000000000";
wait for 1 ns;
clk <= '1';
wait for 1 ns;
clk <= '0';
inA<="000000000000000000000000010000010011100000000000";
inB<="000000000000000000000000010000011010100000000000";
while output_valid = '0' loop
            wait for 1 ns;
            clk <= '1';
            wait for 1 ns;
            clk <= '0';
        end loop;
        for i in 0 to 16384 loop
        wait for 1 ns;
            clk <= '1';
            wait for 1 ns;
            clk <= '0';
        end loop;
        wait;
    end process;
end test;
